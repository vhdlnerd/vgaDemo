library ieee;    use ieee.std_logic_1164.all;


package font_pack is
  -- Define a constant which describes a font table for 256 8x12 characters (and one
  -- for 128 8x16 characters).
  -- Use this later to create a ROM.
  -- For the first font table, all 256 char are defined; so, 12*256=3072 bytes are needed,
  -- but we will round up to the next power of two (4096).  So, other fonts can be defined
  -- here up to 8x16 pixel (all 256 characters).
  -- Note: In Xilinx FPGAs, a 4096 byte ROM will need one or two BRAMs.  Two BRAMs for FPGAs
  --       that only have 18k bit BRAMS -- like the Spartan 3 series.  One BRAM for FPGAs
  --       that have the 36k bit BRAMs -- Virtex 5 and up.
  
  constant FONT_ROM_SIZE : natural := 4096;
  type FontRom_type is array (0 to FONT_ROM_SIZE-1) of std_logic_vector(7 downto 0);
  type Font_type is record
    ID       : natural;
    Width    : natural;
    Height   : natural;
    NumChars : natural;
    Data     : FontRom_type;
  end record Font_type;
 
  constant FONT_ROM_8X12X256 : FontRom_type := (
      -- Char Code: 0x00
    "01111110",  -- 0:  ****** 
    "11000011",  -- 1: **    **
    "10011001",  -- 2: *  **  *
    "10011001",  -- 3: *  **  *
    "11110011",  -- 4: ****  **
    "11100111",  -- 5: ***  ***
    "11100111",  -- 6: ***  ***
    "11111111",  -- 7: ********
    "11100111",  -- 8: ***  ***
    "11100111",  -- 9: ***  ***
    "01111110",  -- A:  ****** 
    "00000000",  -- B:         
      -- Char Code: 0x01
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01110110",  -- 3:  *** ** 
    "11011100",  -- 4: ** ***  
    "00000000",  -- 5:         
    "01110110",  -- 6:  *** ** 
    "11011100",  -- 7: ** ***  
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x02
    "01101110",  -- 0:  ** *** 
    "11011000",  -- 1: ** **   
    "11011000",  -- 2: ** **   
    "11011000",  -- 3: ** **   
    "11011000",  -- 4: ** **   
    "11011110",  -- 5: ** **** 
    "11011000",  -- 6: ** **   
    "11011000",  -- 7: ** **   
    "11011000",  -- 8: ** **   
    "01101110",  -- 9:  ** *** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x03
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01101110",  -- 3:  ** *** 
    "11011011",  -- 4: ** ** **
    "11011011",  -- 5: ** ** **
    "11011111",  -- 6: ** *****
    "11011000",  -- 7: ** **   
    "11011011",  -- 8: ** ** **
    "01101110",  -- 9:  ** *** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x04
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00111000",  -- 3:   ***   
    "01111100",  -- 4:  *****  
    "11111110",  -- 5: ******* 
    "01111100",  -- 6:  *****  
    "00111000",  -- 7:   ***   
    "00010000",  -- 8:    *    
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x05
    "10001000",  -- 0: *   *   
    "10001000",  -- 1: *   *   
    "11111000",  -- 2: *****   
    "10001000",  -- 3: *   *   
    "10001000",  -- 4: *   *   
    "00000000",  -- 5:         
    "00111110",  -- 6:   ***** 
    "00001000",  -- 7:     *   
    "00001000",  -- 8:     *   
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00000000",  -- B:         
      -- Char Code: 0x06
    "11111000",  -- 0: *****   
    "10000000",  -- 1: *       
    "11100000",  -- 2: ***     
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "00000000",  -- 5:         
    "00111110",  -- 6:   ***** 
    "00100000",  -- 7:   *     
    "00111000",  -- 8:   ***   
    "00100000",  -- 9:   *     
    "00100000",  -- A:   *     
    "00000000",  -- B:         
      -- Char Code: 0x07
    "01111000",  -- 0:  ****   
    "10000000",  -- 1: *       
    "10000000",  -- 2: *       
    "10000000",  -- 3: *       
    "01111000",  -- 4:  ****   
    "00000000",  -- 5:         
    "00111100",  -- 6:   ****  
    "00100010",  -- 7:   *   * 
    "00111110",  -- 8:   ***** 
    "00100100",  -- 9:   *  *  
    "00100010",  -- A:   *   * 
    "00000000",  -- B:         
      -- Char Code: 0x08
    "10000000",  -- 0: *       
    "10000000",  -- 1: *       
    "10000000",  -- 2: *       
    "10000000",  -- 3: *       
    "11111000",  -- 4: *****   
    "00000000",  -- 5:         
    "00111110",  -- 6:   ***** 
    "00100000",  -- 7:   *     
    "00111000",  -- 8:   ***   
    "00100000",  -- 9:   *     
    "00100000",  -- A:   *     
    "00000000",  -- B:         
      -- Char Code: 0x09
    "00100010",  -- 0:   *   * 
    "10001000",  -- 1: *   *   
    "00100010",  -- 2:   *   * 
    "10001000",  -- 3: *   *   
    "00100010",  -- 4:   *   * 
    "10001000",  -- 5: *   *   
    "00100010",  -- 6:   *   * 
    "10001000",  -- 7: *   *   
    "00100010",  -- 8:   *   * 
    "10001000",  -- 9: *   *   
    "00100010",  -- A:   *   * 
    "10001000",  -- B: *   *   
      -- Char Code: 0x0A
    "01010101",  -- 0:  * * * *
    "10101010",  -- 1: * * * * 
    "01010101",  -- 2:  * * * *
    "10101010",  -- 3: * * * * 
    "01010101",  -- 4:  * * * *
    "10101010",  -- 5: * * * * 
    "01010101",  -- 6:  * * * *
    "10101010",  -- 7: * * * * 
    "01010101",  -- 8:  * * * *
    "10101010",  -- 9: * * * * 
    "01010101",  -- A:  * * * *
    "10101010",  -- B: * * * * 
      -- Char Code: 0x0B
    "11101110",  -- 0: *** *** 
    "10111011",  -- 1: * *** **
    "11101110",  -- 2: *** *** 
    "10111011",  -- 3: * *** **
    "11101110",  -- 4: *** *** 
    "10111011",  -- 5: * *** **
    "11101110",  -- 6: *** *** 
    "10111011",  -- 7: * *** **
    "11101110",  -- 8: *** *** 
    "10111011",  -- 9: * *** **
    "11101110",  -- A: *** *** 
    "10111011",  -- B: * *** **
      -- Char Code: 0x0C
    "11111111",  -- 0: ********
    "11111111",  -- 1: ********
    "11111111",  -- 2: ********
    "11111111",  -- 3: ********
    "11111111",  -- 4: ********
    "11111111",  -- 5: ********
    "11111111",  -- 6: ********
    "11111111",  -- 7: ********
    "11111111",  -- 8: ********
    "11111111",  -- 9: ********
    "11111111",  -- A: ********
    "11111111",  -- B: ********
      -- Char Code: 0x0D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "11111111",  -- 6: ********
    "11111111",  -- 7: ********
    "11111111",  -- 8: ********
    "11111111",  -- 9: ********
    "11111111",  -- A: ********
    "11111111",  -- B: ********
      -- Char Code: 0x0E
    "11111111",  -- 0: ********
    "11111111",  -- 1: ********
    "11111111",  -- 2: ********
    "11111111",  -- 3: ********
    "11111111",  -- 4: ********
    "11111111",  -- 5: ********
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x0F
    "11110000",  -- 0: ****    
    "11110000",  -- 1: ****    
    "11110000",  -- 2: ****    
    "11110000",  -- 3: ****    
    "11110000",  -- 4: ****    
    "11110000",  -- 5: ****    
    "11110000",  -- 6: ****    
    "11110000",  -- 7: ****    
    "11110000",  -- 8: ****    
    "11110000",  -- 9: ****    
    "11110000",  -- A: ****    
    "11110000",  -- B: ****    
      -- Char Code: 0x10
    "00001111",  -- 0:     ****
    "00001111",  -- 1:     ****
    "00001111",  -- 2:     ****
    "00001111",  -- 3:     ****
    "00001111",  -- 4:     ****
    "00001111",  -- 5:     ****
    "00001111",  -- 6:     ****
    "00001111",  -- 7:     ****
    "00001111",  -- 8:     ****
    "00001111",  -- 9:     ****
    "00001111",  -- A:     ****
    "00001111",  -- B:     ****
      -- Char Code: 0x11
    "10001000",  -- 0: *   *   
    "11001000",  -- 1: **  *   
    "10101000",  -- 2: * * *   
    "10011000",  -- 3: *  **   
    "10001000",  -- 4: *   *   
    "00000000",  -- 5:         
    "00100000",  -- 6:   *     
    "00100000",  -- 7:   *     
    "00100000",  -- 8:   *     
    "00100000",  -- 9:   *     
    "00111110",  -- A:   ***** 
    "00000000",  -- B:         
      -- Char Code: 0x12
    "10001000",  -- 0: *   *   
    "10001000",  -- 1: *   *   
    "01010000",  -- 2:  * *    
    "01010000",  -- 3:  * *    
    "00100000",  -- 4:   *     
    "00000000",  -- 5:         
    "00111110",  -- 6:   ***** 
    "00001000",  -- 7:     *   
    "00001000",  -- 8:     *   
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00000000",  -- B:         
      -- Char Code: 0x13
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000110",  -- 2:      ** 
    "00001100",  -- 3:     **  
    "00011000",  -- 4:    **   
    "00110000",  -- 5:   **    
    "01111110",  -- 6:  ****** 
    "00000000",  -- 7:         
    "01111110",  -- 8:  ****** 
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x14
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01100000",  -- 2:  **     
    "00110000",  -- 3:   **    
    "00011000",  -- 4:    **   
    "00001100",  -- 5:     **  
    "01111110",  -- 6:  ****** 
    "00000000",  -- 7:         
    "01111110",  -- 8:  ****** 
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x15
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000110",  -- 2:      ** 
    "00001100",  -- 3:     **  
    "11111110",  -- 4: ******* 
    "00111000",  -- 5:   ***   
    "11111110",  -- 6: ******* 
    "01100000",  -- 7:  **     
    "11000000",  -- 8: **      
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x16
    "00000000",  -- 0:         
    "00000010",  -- 1:       * 
    "00001110",  -- 2:     *** 
    "00111110",  -- 3:   ***** 
    "01111110",  -- 4:  ****** 
    "11111110",  -- 5: ******* 
    "01111110",  -- 6:  ****** 
    "00111110",  -- 7:   ***** 
    "00001110",  -- 8:     *** 
    "00000010",  -- 9:       * 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x17
    "00000000",  -- 0:         
    "10000000",  -- 1: *       
    "11100000",  -- 2: ***     
    "11110000",  -- 3: ****    
    "11111100",  -- 4: ******  
    "11111110",  -- 5: ******* 
    "11111100",  -- 6: ******  
    "11110000",  -- 7: ****    
    "11100000",  -- 8: ***     
    "10000000",  -- 9: *       
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x18
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00111100",  -- 2:   ****  
    "01111110",  -- 3:  ****** 
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x19
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "01111110",  -- 7:  ****** 
    "00111100",  -- 8:   ****  
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x1A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00011000",  -- 3:    **   
    "00001100",  -- 4:     **  
    "11111110",  -- 5: ******* 
    "00001100",  -- 6:     **  
    "00011000",  -- 7:    **   
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x1B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00110000",  -- 3:   **    
    "01100000",  -- 4:  **     
    "11111110",  -- 5: ******* 
    "01100000",  -- 6:  **     
    "00110000",  -- 7:   **    
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x1C
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00111100",  -- 2:   ****  
    "01111110",  -- 3:  ****** 
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "01111110",  -- 7:  ****** 
    "00111100",  -- 8:   ****  
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x1D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00101000",  -- 3:   * *   
    "01101100",  -- 4:  ** **  
    "11111110",  -- 5: ******* 
    "01101100",  -- 6:  ** **  
    "00101000",  -- 7:   * *   
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x1E
    "00000000",  -- 0:         
    "00000110",  -- 1:      ** 
    "00000110",  -- 2:      ** 
    "00110110",  -- 3:   ** ** 
    "01100110",  -- 4:  **  ** 
    "11111110",  -- 5: ******* 
    "01100000",  -- 6:  **     
    "00110000",  -- 7:   **    
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x1F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "11000000",  -- 3: **      
    "01111100",  -- 4:  *****  
    "01101110",  -- 5:  ** *** 
    "01101100",  -- 6:  ** **  
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x20
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x21
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00111100",  -- 2:   ****  
    "00111100",  -- 3:   ****  
    "00111100",  -- 4:   ****  
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00000000",  -- 7:         
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x22
    "00000000",  -- 0:         
    "00110110",  -- 1:   ** ** 
    "00110110",  -- 2:   ** ** 
    "00010100",  -- 3:    * *  
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x23
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01101100",  -- 3:  ** **  
    "11111110",  -- 4: ******* 
    "01101100",  -- 5:  ** **  
    "01101100",  -- 6:  ** **  
    "01101100",  -- 7:  ** **  
    "11111110",  -- 8: ******* 
    "01101100",  -- 9:  ** **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x24
    "00000000",  -- 0:         
    "00010000",  -- 1:    *    
    "01111100",  -- 2:  *****  
    "11010110",  -- 3: ** * ** 
    "01110000",  -- 4:  ***    
    "00111000",  -- 5:   ***   
    "00011100",  -- 6:    ***  
    "11010110",  -- 7: ** * ** 
    "01111100",  -- 8:  *****  
    "00010000",  -- 9:    *    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x25
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01100010",  -- 3:  **   * 
    "01100110",  -- 4:  **  ** 
    "00001100",  -- 5:     **  
    "00011000",  -- 6:    **   
    "00110000",  -- 7:   **    
    "01100110",  -- 8:  **  ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x26
    "00000000",  -- 0:         
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "00111000",  -- 3:   ***   
    "00111000",  -- 4:   ***   
    "01110010",  -- 5:  ***  * 
    "11111110",  -- 6: ******* 
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x27
    "00011100",  -- 0:    ***  
    "00011100",  -- 1:    ***  
    "00001100",  -- 2:     **  
    "00011000",  -- 3:    **   
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x28
    "00000000",  -- 0:         
    "00001100",  -- 1:     **  
    "00011000",  -- 2:    **   
    "00110000",  -- 3:   **    
    "00110000",  -- 4:   **    
    "00110000",  -- 5:   **    
    "00110000",  -- 6:   **    
    "00110000",  -- 7:   **    
    "00011000",  -- 8:    **   
    "00001100",  -- 9:     **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x29
    "00000000",  -- 0:         
    "00110000",  -- 1:   **    
    "00011000",  -- 2:    **   
    "00001100",  -- 3:     **  
    "00001100",  -- 4:     **  
    "00001100",  -- 5:     **  
    "00001100",  -- 6:     **  
    "00001100",  -- 7:     **  
    "00011000",  -- 8:    **   
    "00110000",  -- 9:   **    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x2A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01101100",  -- 3:  ** **  
    "00111000",  -- 4:   ***   
    "11111110",  -- 5: ******* 
    "00111000",  -- 6:   ***   
    "01101100",  -- 7:  ** **  
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x2B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "01111110",  -- 5:  ****** 
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x2C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00001100",  -- 7:     **  
    "00001100",  -- 8:     **  
    "00001100",  -- 9:     **  
    "00011000",  -- A:    **   
    "00000000",  -- B:         
      -- Char Code: 0x2D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "11111110",  -- 5: ******* 
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x2E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x2F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000110",  -- 3:      ** 
    "00001100",  -- 4:     **  
    "00011000",  -- 5:    **   
    "00110000",  -- 6:   **    
    "01100000",  -- 7:  **     
    "11000000",  -- 8: **      
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x30
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11010110",  -- 5: ** * ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x31
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "01111000",  -- 2:  ****   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x32
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "00001100",  -- 4:     **  
    "00011000",  -- 5:    **   
    "00110000",  -- 6:   **    
    "01100000",  -- 7:  **     
    "11000110",  -- 8: **   ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x33
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "00000110",  -- 3:      ** 
    "00000110",  -- 4:      ** 
    "00111100",  -- 5:   ****  
    "00000110",  -- 6:      ** 
    "00000110",  -- 7:      ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x34
    "00000000",  -- 0:         
    "00001100",  -- 1:     **  
    "00011100",  -- 2:    ***  
    "00111100",  -- 3:   ****  
    "01101100",  -- 4:  ** **  
    "11001100",  -- 5: **  **  
    "11111110",  -- 6: ******* 
    "00001100",  -- 7:     **  
    "00001100",  -- 8:     **  
    "00001100",  -- 9:     **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x35
    "00000000",  -- 0:         
    "11111110",  -- 1: ******* 
    "11000000",  -- 2: **      
    "11000000",  -- 3: **      
    "11000000",  -- 4: **      
    "11111100",  -- 5: ******  
    "00000110",  -- 6:      ** 
    "00000110",  -- 7:      ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x36
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000000",  -- 3: **      
    "11000000",  -- 4: **      
    "11111100",  -- 5: ******  
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x37
    "00000000",  -- 0:         
    "11111110",  -- 1: ******* 
    "11000110",  -- 2: **   ** 
    "00001100",  -- 3:     **  
    "00011000",  -- 4:    **   
    "00110000",  -- 5:   **    
    "00110000",  -- 6:   **    
    "00110000",  -- 7:   **    
    "00110000",  -- 8:   **    
    "00110000",  -- 9:   **    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x38
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "01111100",  -- 5:  *****  
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x39
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "01111110",  -- 5:  ****** 
    "00000110",  -- 6:      ** 
    "00000110",  -- 7:      ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x3A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00001100",  -- 3:     **  
    "00001100",  -- 4:     **  
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00001100",  -- 7:     **  
    "00001100",  -- 8:     **  
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x3B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00001100",  -- 3:     **  
    "00001100",  -- 4:     **  
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00001100",  -- 7:     **  
    "00001100",  -- 8:     **  
    "00001100",  -- 9:     **  
    "00011000",  -- A:    **   
    "00000000",  -- B:         
      -- Char Code: 0x3C
    "00000000",  -- 0:         
    "00001100",  -- 1:     **  
    "00011000",  -- 2:    **   
    "00110000",  -- 3:   **    
    "01100000",  -- 4:  **     
    "11000000",  -- 5: **      
    "01100000",  -- 6:  **     
    "00110000",  -- 7:   **    
    "00011000",  -- 8:    **   
    "00001100",  -- 9:     **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x3D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111110",  -- 4: ******* 
    "00000000",  -- 5:         
    "11111110",  -- 6: ******* 
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x3E
    "00000000",  -- 0:         
    "01100000",  -- 1:  **     
    "00110000",  -- 2:   **    
    "00011000",  -- 3:    **   
    "00001100",  -- 4:     **  
    "00000110",  -- 5:      ** 
    "00001100",  -- 6:     **  
    "00011000",  -- 7:    **   
    "00110000",  -- 8:   **    
    "01100000",  -- 9:  **     
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x3F
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "00001100",  -- 4:     **  
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00000000",  -- 7:         
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x40
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11011110",  -- 4: ** **** 
    "11011110",  -- 5: ** **** 
    "11011110",  -- 6: ** **** 
    "11011100",  -- 7: ** ***  
    "11000000",  -- 8: **      
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x41
    "00000000",  -- 0:         
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11111110",  -- 6: ******* 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x42
    "00000000",  -- 0:         
    "11111100",  -- 1: ******  
    "01100110",  -- 2:  **  ** 
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01111100",  -- 5:  *****  
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01100110",  -- 8:  **  ** 
    "11111100",  -- 9: ******  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x43
    "00000000",  -- 0:         
    "00111100",  -- 1:   ****  
    "01100110",  -- 2:  **  ** 
    "11000000",  -- 3: **      
    "11000000",  -- 4: **      
    "11000000",  -- 5: **      
    "11000000",  -- 6: **      
    "11000000",  -- 7: **      
    "01100110",  -- 8:  **  ** 
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x44
    "00000000",  -- 0:         
    "11111000",  -- 1: *****   
    "01101100",  -- 2:  ** **  
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01101100",  -- 8:  ** **  
    "11111000",  -- 9: *****   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x45
    "00000000",  -- 0:         
    "11111110",  -- 1: ******* 
    "01100110",  -- 2:  **  ** 
    "01100000",  -- 3:  **     
    "01100000",  -- 4:  **     
    "01111100",  -- 5:  *****  
    "01100000",  -- 6:  **     
    "01100000",  -- 7:  **     
    "01100110",  -- 8:  **  ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x46
    "00000000",  -- 0:         
    "11111110",  -- 1: ******* 
    "01100110",  -- 2:  **  ** 
    "01100000",  -- 3:  **     
    "01100000",  -- 4:  **     
    "01111100",  -- 5:  *****  
    "01100000",  -- 6:  **     
    "01100000",  -- 7:  **     
    "01100000",  -- 8:  **     
    "11110000",  -- 9: ****    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x47
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000000",  -- 4: **      
    "11000000",  -- 5: **      
    "11001110",  -- 6: **  *** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x48
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11111110",  -- 5: ******* 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x49
    "00000000",  -- 0:         
    "00111100",  -- 1:   ****  
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x4A
    "00000000",  -- 0:         
    "00111100",  -- 1:   ****  
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "11011000",  -- 7: ** **   
    "11011000",  -- 8: ** **   
    "01110000",  -- 9:  ***    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x4B
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11001100",  -- 2: **  **  
    "11011000",  -- 3: ** **   
    "11110000",  -- 4: ****    
    "11110000",  -- 5: ****    
    "11011000",  -- 6: ** **   
    "11001100",  -- 7: **  **  
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x4C
    "00000000",  -- 0:         
    "11110000",  -- 1: ****    
    "01100000",  -- 2:  **     
    "01100000",  -- 3:  **     
    "01100000",  -- 4:  **     
    "01100000",  -- 5:  **     
    "01100000",  -- 6:  **     
    "01100010",  -- 7:  **   * 
    "01100110",  -- 8:  **  ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x4D
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "11101110",  -- 3: *** *** 
    "11111110",  -- 4: ******* 
    "11010110",  -- 5: ** * ** 
    "11010110",  -- 6: ** * ** 
    "11010110",  -- 7: ** * ** 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x4E
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "11100110",  -- 3: ***  ** 
    "11100110",  -- 4: ***  ** 
    "11110110",  -- 5: **** ** 
    "11011110",  -- 6: ** **** 
    "11001110",  -- 7: **  *** 
    "11001110",  -- 8: **  *** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x4F
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x50
    "00000000",  -- 0:         
    "11111100",  -- 1: ******  
    "01100110",  -- 2:  **  ** 
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01111100",  -- 5:  *****  
    "01100000",  -- 6:  **     
    "01100000",  -- 7:  **     
    "01100000",  -- 8:  **     
    "11110000",  -- 9: ****    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x51
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11010110",  -- 8: ** * ** 
    "01111100",  -- 9:  *****  
    "00000110",  -- A:      ** 
    "00000000",  -- B:         
      -- Char Code: 0x52
    "00000000",  -- 0:         
    "11111100",  -- 1: ******  
    "01100110",  -- 2:  **  ** 
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01111100",  -- 5:  *****  
    "01111000",  -- 6:  ****   
    "01101100",  -- 7:  ** **  
    "01100110",  -- 8:  **  ** 
    "11100110",  -- 9: ***  ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x53
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000000",  -- 3: **      
    "01100000",  -- 4:  **     
    "00111000",  -- 5:   ***   
    "00001100",  -- 6:     **  
    "00000110",  -- 7:      ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x54
    "00000000",  -- 0:         
    "01111110",  -- 1:  ****** 
    "01011010",  -- 2:  * ** * 
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x55
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x56
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "01101100",  -- 7:  ** **  
    "00111000",  -- 8:   ***   
    "00010000",  -- 9:    *    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x57
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "11010110",  -- 3: ** * ** 
    "11010110",  -- 4: ** * ** 
    "11010110",  -- 5: ** * ** 
    "11111110",  -- 6: ******* 
    "11101110",  -- 7: *** *** 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x58
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "01101100",  -- 3:  ** **  
    "00111000",  -- 4:   ***   
    "00111000",  -- 5:   ***   
    "00111000",  -- 6:   ***   
    "01101100",  -- 7:  ** **  
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x59
    "00000000",  -- 0:         
    "01100110",  -- 1:  **  ** 
    "01100110",  -- 2:  **  ** 
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "00111100",  -- 5:   ****  
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x5A
    "00000000",  -- 0:         
    "11111110",  -- 1: ******* 
    "11000110",  -- 2: **   ** 
    "10001100",  -- 3: *   **  
    "00011000",  -- 4:    **   
    "00110000",  -- 5:   **    
    "01100000",  -- 6:  **     
    "11000010",  -- 7: **    * 
    "11000110",  -- 8: **   ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x5B
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "01100000",  -- 2:  **     
    "01100000",  -- 3:  **     
    "01100000",  -- 4:  **     
    "01100000",  -- 5:  **     
    "01100000",  -- 6:  **     
    "01100000",  -- 7:  **     
    "01100000",  -- 8:  **     
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x5C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "11000000",  -- 3: **      
    "01100000",  -- 4:  **     
    "00110000",  -- 5:   **    
    "00011000",  -- 6:    **   
    "00001100",  -- 7:     **  
    "00000110",  -- 8:      ** 
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x5D
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "00001100",  -- 2:     **  
    "00001100",  -- 3:     **  
    "00001100",  -- 4:     **  
    "00001100",  -- 5:     **  
    "00001100",  -- 6:     **  
    "00001100",  -- 7:     **  
    "00001100",  -- 8:     **  
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x5E
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00111100",  -- 2:   ****  
    "01100110",  -- 3:  **  ** 
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x5F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "11111111",  -- B: ********
      -- Char Code: 0x60
    "00011100",  -- 0:    ***  
    "00011100",  -- 1:    ***  
    "00011000",  -- 2:    **   
    "00001100",  -- 3:     **  
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x61
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x62
    "00000000",  -- 0:         
    "11100000",  -- 1: ***     
    "01100000",  -- 2:  **     
    "01100000",  -- 3:  **     
    "01111100",  -- 4:  *****  
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01100110",  -- 8:  **  ** 
    "11111100",  -- 9: ******  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x63
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000000",  -- 6: **      
    "11000000",  -- 7: **      
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x64
    "00000000",  -- 0:         
    "00011100",  -- 1:    ***  
    "00001100",  -- 2:     **  
    "00001100",  -- 3:     **  
    "01111100",  -- 4:  *****  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x65
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11111110",  -- 6: ******* 
    "11000000",  -- 7: **      
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x66
    "00000000",  -- 0:         
    "00011100",  -- 1:    ***  
    "00110110",  -- 2:   ** ** 
    "00110000",  -- 3:   **    
    "00110000",  -- 4:   **    
    "11111100",  -- 5: ******  
    "00110000",  -- 6:   **    
    "00110000",  -- 7:   **    
    "00110000",  -- 8:   **    
    "01111000",  -- 9:  ****   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x67
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01110110",  -- 4:  *** ** 
    "11001110",  -- 5: **  *** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "01111110",  -- 8:  ****** 
    "00000110",  -- 9:      ** 
    "11000110",  -- A: **   ** 
    "01111100",  -- B:  *****  
      -- Char Code: 0x68
    "00000000",  -- 0:         
    "11100000",  -- 1: ***     
    "01100000",  -- 2:  **     
    "01100000",  -- 3:  **     
    "01101100",  -- 4:  ** **  
    "01110110",  -- 5:  *** ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01100110",  -- 8:  **  ** 
    "11100110",  -- 9: ***  ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x69
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00000000",  -- 3:         
    "00111000",  -- 4:   ***   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x6A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00001100",  -- 2:     **  
    "00001100",  -- 3:     **  
    "00000000",  -- 4:         
    "00011100",  -- 5:    ***  
    "00001100",  -- 6:     **  
    "00001100",  -- 7:     **  
    "00001100",  -- 8:     **  
    "11001100",  -- 9: **  **  
    "11001100",  -- A: **  **  
    "01111000",  -- B:  ****   
      -- Char Code: 0x6B
    "00000000",  -- 0:         
    "11100000",  -- 1: ***     
    "01100000",  -- 2:  **     
    "01100000",  -- 3:  **     
    "01100110",  -- 4:  **  ** 
    "01101100",  -- 5:  ** **  
    "01111000",  -- 6:  ****   
    "01101100",  -- 7:  ** **  
    "01100110",  -- 8:  **  ** 
    "11100110",  -- 9: ***  ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x6C
    "00000000",  -- 0:         
    "01110000",  -- 1:  ***    
    "00110000",  -- 2:   **    
    "00110000",  -- 3:   **    
    "00110000",  -- 4:   **    
    "00110000",  -- 5:   **    
    "00110000",  -- 6:   **    
    "00110000",  -- 7:   **    
    "00110100",  -- 8:   ** *  
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x6D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01101100",  -- 4:  ** **  
    "11111110",  -- 5: ******* 
    "11010110",  -- 6: ** * ** 
    "11010110",  -- 7: ** * ** 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x6E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11011100",  -- 4: ** ***  
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01100110",  -- 8:  **  ** 
    "01100110",  -- 9:  **  ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x6F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x70
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11011100",  -- 4: ** ***  
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01111100",  -- 8:  *****  
    "01100000",  -- 9:  **     
    "01100000",  -- A:  **     
    "11110000",  -- B: ****    
      -- Char Code: 0x71
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01110110",  -- 4:  *** ** 
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "01111100",  -- 8:  *****  
    "00001100",  -- 9:     **  
    "00001100",  -- A:     **  
    "00011110",  -- B:    **** 
      -- Char Code: 0x72
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11011100",  -- 4: ** ***  
    "01100110",  -- 5:  **  ** 
    "01100000",  -- 6:  **     
    "01100000",  -- 7:  **     
    "01100000",  -- 8:  **     
    "11110000",  -- 9: ****    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x73
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "01110000",  -- 6:  ***    
    "00011100",  -- 7:    ***  
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x74
    "00000000",  -- 0:         
    "00110000",  -- 1:   **    
    "00110000",  -- 2:   **    
    "00110000",  -- 3:   **    
    "11111100",  -- 4: ******  
    "00110000",  -- 5:   **    
    "00110000",  -- 6:   **    
    "00110000",  -- 7:   **    
    "00110110",  -- 8:   ** ** 
    "00011100",  -- 9:    ***  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x75
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11001100",  -- 4: **  **  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x76
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "01101100",  -- 7:  ** **  
    "00111000",  -- 8:   ***   
    "00010000",  -- 9:    *    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x77
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11010110",  -- 6: ** * ** 
    "11010110",  -- 7: ** * ** 
    "11111110",  -- 8: ******* 
    "01101100",  -- 9:  ** **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x78
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11000110",  -- 4: **   ** 
    "01101100",  -- 5:  ** **  
    "00111000",  -- 6:   ***   
    "00111000",  -- 7:   ***   
    "01101100",  -- 8:  ** **  
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x79
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11001110",  -- 7: **  *** 
    "01110110",  -- 8:  *** ** 
    "00000110",  -- 9:      ** 
    "11000110",  -- A: **   ** 
    "01111100",  -- B:  *****  
      -- Char Code: 0x7A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111110",  -- 4: ******* 
    "10001100",  -- 5: *   **  
    "00011000",  -- 6:    **   
    "00110000",  -- 7:   **    
    "01100010",  -- 8:  **   * 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x7B
    "00000000",  -- 0:         
    "00001110",  -- 1:     *** 
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "01110000",  -- 5:  ***    
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00001110",  -- 9:     *** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x7C
    "00000000",  -- 0:         
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x7D
    "00000000",  -- 0:         
    "01110000",  -- 1:  ***    
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00001110",  -- 5:     *** 
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "01110000",  -- 9:  ***    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x7E
    "00000000",  -- 0:         
    "01110110",  -- 1:  *** ** 
    "11011100",  -- 2: ** ***  
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x7F
    "01100110",  -- 0:  **  ** 
    "01100110",  -- 1:  **  ** 
    "00000000",  -- 2:         
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01100110",  -- 5:  **  ** 
    "00111100",  -- 6:   ****  
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x80
    "00110000",  -- 0:   **    
    "00011000",  -- 1:    **   
    "00000000",  -- 2:         
    "00111000",  -- 3:   ***   
    "01101100",  -- 4:  ** **  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11111110",  -- 7: ******* 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x81
    "00011000",  -- 0:    **   
    "00110000",  -- 1:   **    
    "00000000",  -- 2:         
    "00111000",  -- 3:   ***   
    "01101100",  -- 4:  ** **  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11111110",  -- 7: ******* 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x82
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "00111000",  -- 2:   ***   
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11111110",  -- 7: ******* 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x83
    "01110110",  -- 0:  *** ** 
    "11011100",  -- 1: ** ***  
    "00000000",  -- 2:         
    "00111000",  -- 3:   ***   
    "01101100",  -- 4:  ** **  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11111110",  -- 7: ******* 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x84
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "00111000",  -- 3:   ***   
    "01101100",  -- 4:  ** **  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11111110",  -- 7: ******* 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x85
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "00111000",  -- 2:   ***   
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11111110",  -- 7: ******* 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x86
    "01111110",  -- 0:  ****** 
    "11011000",  -- 1: ** **   
    "11011000",  -- 2: ** **   
    "11011000",  -- 3: ** **   
    "11011000",  -- 4: ** **   
    "11111110",  -- 5: ******* 
    "11011000",  -- 6: ** **   
    "11011000",  -- 7: ** **   
    "11011000",  -- 8: ** **   
    "11011110",  -- 9: ** **** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x87
    "00000000",  -- 0:         
    "00111100",  -- 1:   ****  
    "01100110",  -- 2:  **  ** 
    "11000000",  -- 3: **      
    "11000000",  -- 4: **      
    "11000000",  -- 5: **      
    "11000110",  -- 6: **   ** 
    "01100110",  -- 7:  **  ** 
    "00111100",  -- 8:   ****  
    "00011000",  -- 9:    **   
    "11001100",  -- A: **  **  
    "00111000",  -- B:   ***   
      -- Char Code: 0x88
    "00011000",  -- 0:    **   
    "00001100",  -- 1:     **  
    "00000000",  -- 2:         
    "11111110",  -- 3: ******* 
    "01100110",  -- 4:  **  ** 
    "01100000",  -- 5:  **     
    "01111100",  -- 6:  *****  
    "01100000",  -- 7:  **     
    "01100110",  -- 8:  **  ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x89
    "00011000",  -- 0:    **   
    "00110000",  -- 1:   **    
    "00000000",  -- 2:         
    "11111110",  -- 3: ******* 
    "01100110",  -- 4:  **  ** 
    "01100000",  -- 5:  **     
    "01111100",  -- 6:  *****  
    "01100000",  -- 7:  **     
    "01100110",  -- 8:  **  ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x8A
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "11111110",  -- 3: ******* 
    "01100110",  -- 4:  **  ** 
    "01100000",  -- 5:  **     
    "01111100",  -- 6:  *****  
    "01100000",  -- 7:  **     
    "01100110",  -- 8:  **  ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x8B
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "11111110",  -- 3: ******* 
    "01100110",  -- 4:  **  ** 
    "01100000",  -- 5:  **     
    "01111100",  -- 6:  *****  
    "01100000",  -- 7:  **     
    "01100110",  -- 8:  **  ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x8C
    "00011000",  -- 0:    **   
    "00001100",  -- 1:     **  
    "00000000",  -- 2:         
    "00111100",  -- 3:   ****  
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x8D
    "00011000",  -- 0:    **   
    "00110000",  -- 1:   **    
    "00000000",  -- 2:         
    "00111100",  -- 3:   ****  
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x8E
    "00111100",  -- 0:   ****  
    "01100110",  -- 1:  **  ** 
    "00000000",  -- 2:         
    "00111100",  -- 3:   ****  
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x8F
    "01100110",  -- 0:  **  ** 
    "01100110",  -- 1:  **  ** 
    "00000000",  -- 2:         
    "00111100",  -- 3:   ****  
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x90
    "00000000",  -- 0:         
    "11111000",  -- 1: *****   
    "01101100",  -- 2:  ** **  
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "11110110",  -- 5: **** ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01101100",  -- 8:  ** **  
    "11111000",  -- 9: *****   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x91
    "01110110",  -- 0:  *** ** 
    "11011100",  -- 1: ** ***  
    "00000000",  -- 2:         
    "11000110",  -- 3: **   ** 
    "11100110",  -- 4: ***  ** 
    "11110110",  -- 5: **** ** 
    "11011110",  -- 6: ** **** 
    "11001110",  -- 7: **  *** 
    "11000110",  -- 8: **   ** 
    "11000110",  -- 9: **   ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x92
    "00110000",  -- 0:   **    
    "00011000",  -- 1:    **   
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x93
    "00011000",  -- 0:    **   
    "00110000",  -- 1:   **    
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x94
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x95
    "01110110",  -- 0:  *** ** 
    "11011100",  -- 1: ** ***  
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x96
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x97
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01101100",  -- 4:  ** **  
    "00111000",  -- 5:   ***   
    "00111000",  -- 6:   ***   
    "01101100",  -- 7:  ** **  
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x98
    "00000000",  -- 0:         
    "01111110",  -- 1:  ****** 
    "11000110",  -- 2: **   ** 
    "11001110",  -- 3: **  *** 
    "11011110",  -- 4: ** **** 
    "11010110",  -- 5: ** * ** 
    "11110110",  -- 6: **** ** 
    "11100110",  -- 7: ***  ** 
    "11000110",  -- 8: **   ** 
    "11111100",  -- 9: ******  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x99
    "00110000",  -- 0:   **    
    "00011000",  -- 1:    **   
    "00000000",  -- 2:         
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x9A
    "00011000",  -- 0:    **   
    "00110000",  -- 1:   **    
    "00000000",  -- 2:         
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x9B
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x9C
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "00000000",  -- 2:         
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x9D
    "00001100",  -- 0:     **  
    "00011000",  -- 1:    **   
    "00000000",  -- 2:         
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01100110",  -- 5:  **  ** 
    "00111100",  -- 6:   ****  
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x9E
    "00000000",  -- 0:         
    "11110000",  -- 1: ****    
    "01100000",  -- 2:  **     
    "01111100",  -- 3:  *****  
    "01100110",  -- 4:  **  ** 
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "01111100",  -- 7:  *****  
    "01100000",  -- 8:  **     
    "11110000",  -- 9: ****    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0x9F
    "00000000",  -- 0:         
    "01111100",  -- 1:  *****  
    "11000110",  -- 2: **   ** 
    "11000110",  -- 3: **   ** 
    "11000110",  -- 4: **   ** 
    "11001100",  -- 5: **  **  
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11010110",  -- 8: ** * ** 
    "11011100",  -- 9: ** ***  
    "10000000",  -- A: *       
    "00000000",  -- B:         
      -- Char Code: 0xA0
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "10000010",  -- 9: *     * 
    "11111110",  -- A: ******* 
    "00000000",  -- B:         
      -- Char Code: 0xA1
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00000000",  -- 5:         
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00111100",  -- 8:   ****  
    "00111100",  -- 9:   ****  
    "00111100",  -- A:   ****  
    "00011000",  -- B:    **   
      -- Char Code: 0xA2
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "01111100",  -- 3:  *****  
    "11010110",  -- 4: ** * ** 
    "11010000",  -- 5: ** *    
    "11010000",  -- 6: ** *    
    "11010110",  -- 7: ** * ** 
    "01111100",  -- 8:  *****  
    "00010000",  -- 9:    *    
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xA3
    "00000000",  -- 0:         
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "01100000",  -- 3:  **     
    "01100000",  -- 4:  **     
    "11110000",  -- 5: ****    
    "01100000",  -- 6:  **     
    "01100110",  -- 7:  **  ** 
    "11110110",  -- 8: **** ** 
    "01101100",  -- 9:  ** **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xA4
    "00000000",  -- 0:         
    "00111100",  -- 1:   ****  
    "01100010",  -- 2:  **   * 
    "01100000",  -- 3:  **     
    "11111000",  -- 4: *****   
    "01100000",  -- 5:  **     
    "11111000",  -- 6: *****   
    "01100000",  -- 7:  **     
    "01100010",  -- 8:  **   * 
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xA5
    "00000000",  -- 0:         
    "01100110",  -- 1:  **  ** 
    "01100110",  -- 2:  **  ** 
    "00111100",  -- 3:   ****  
    "00011000",  -- 4:    **   
    "01111110",  -- 5:  ****** 
    "00011000",  -- 6:    **   
    "00111100",  -- 7:   ****  
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xA6
    "01101100",  -- 0:  ** **  
    "00111000",  -- 1:   ***   
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000000",  -- 5: **      
    "01111100",  -- 6:  *****  
    "00000110",  -- 7:      ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xA7
    "01111100",  -- 0:  *****  
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "01100000",  -- 3:  **     
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "01111100",  -- 7:  *****  
    "00001100",  -- 8:     **  
    "11000110",  -- 9: **   ** 
    "11000110",  -- A: **   ** 
    "01111100",  -- B:  *****  
      -- Char Code: 0xA8
    "00000000",  -- 0:         
    "01101100",  -- 1:  ** **  
    "00111000",  -- 2:   ***   
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "01110000",  -- 6:  ***    
    "00011100",  -- 7:    ***  
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xA9
    "01111110",  -- 0:  ****** 
    "10000001",  -- 1: *      *
    "10011001",  -- 2: *  **  *
    "10100101",  -- 3: * *  * *
    "10100001",  -- 4: * *    *
    "10100001",  -- 5: * *    *
    "10100101",  -- 6: * *  * *
    "10011001",  -- 7: *  **  *
    "10000001",  -- 8: *      *
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xAA
    "00111100",  -- 0:   ****  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "00111110",  -- 3:   ***** 
    "00000000",  -- 4:         
    "01111110",  -- 5:  ****** 
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xAB
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00110110",  -- 3:   ** ** 
    "01101100",  -- 4:  ** **  
    "11011000",  -- 5: ** **   
    "01101100",  -- 6:  ** **  
    "00110110",  -- 7:   ** ** 
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xAC
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "01111110",  -- 5:  ****** 
    "00000110",  -- 6:      ** 
    "00000110",  -- 7:      ** 
    "00000110",  -- 8:      ** 
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xAD
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "01111110",  -- 5:  ****** 
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xAE
    "01111110",  -- 0:  ****** 
    "10000001",  -- 1: *      *
    "10111001",  -- 2: * ***  *
    "10100101",  -- 3: * *  * *
    "10100101",  -- 4: * *  * *
    "10111001",  -- 5: * ***  *
    "10100101",  -- 6: * *  * *
    "10100101",  -- 7: * *  * *
    "10000001",  -- 8: *      *
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xAF
    "11111111",  -- 0: ********
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB0
    "00000000",  -- 0:         
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "00111000",  -- 3:   ***   
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB1
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "01111110",  -- 5:  ****** 
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00000000",  -- 8:         
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB2
    "00000000",  -- 0:         
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "00011000",  -- 3:    **   
    "00110000",  -- 4:   **    
    "01111100",  -- 5:  *****  
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB3
    "00000000",  -- 0:         
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "00011000",  -- 3:    **   
    "01101100",  -- 4:  ** **  
    "00111000",  -- 5:   ***   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB4
    "01101100",  -- 0:  ** **  
    "00111000",  -- 1:   ***   
    "00000000",  -- 2:         
    "11111110",  -- 3: ******* 
    "11000110",  -- 4: **   ** 
    "00001100",  -- 5:     **  
    "00111000",  -- 6:   ***   
    "01100010",  -- 7:  **   * 
    "11000110",  -- 8: **   ** 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB5
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11001100",  -- 4: **  **  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "11110110",  -- 9: **** ** 
    "11000000",  -- A: **      
    "11000000",  -- B: **      
      -- Char Code: 0xB6
    "00000000",  -- 0:         
    "01111111",  -- 1:  *******
    "11011011",  -- 2: ** ** **
    "11011011",  -- 3: ** ** **
    "11011011",  -- 4: ** ** **
    "01111011",  -- 5:  **** **
    "00011011",  -- 6:    ** **
    "00011011",  -- 7:    ** **
    "00011011",  -- 8:    ** **
    "00011011",  -- 9:    ** **
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB7
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB8
    "00000000",  -- 0:         
    "01101100",  -- 1:  ** **  
    "00111000",  -- 2:   ***   
    "00000000",  -- 3:         
    "11111110",  -- 4: ******* 
    "10001100",  -- 5: *   **  
    "00011000",  -- 6:    **   
    "00110000",  -- 7:   **    
    "01100010",  -- 8:  **   * 
    "11111110",  -- 9: ******* 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xB9
    "00000000",  -- 0:         
    "00110000",  -- 1:   **    
    "01110000",  -- 2:  ***    
    "00110000",  -- 3:   **    
    "00110000",  -- 4:   **    
    "01111000",  -- 5:  ****   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xBA
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "00111000",  -- 3:   ***   
    "00000000",  -- 4:         
    "01111100",  -- 5:  *****  
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xBB
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "11011000",  -- 3: ** **   
    "01101100",  -- 4:  ** **  
    "00110110",  -- 5:   ** ** 
    "01101100",  -- 6:  ** **  
    "11011000",  -- 7: ** **   
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xBC
    "00000000",  -- 0:         
    "01101110",  -- 1:  ** *** 
    "11011011",  -- 2: ** ** **
    "11011011",  -- 3: ** ** **
    "11011111",  -- 4: ** *****
    "11011000",  -- 5: ** **   
    "11011000",  -- 6: ** **   
    "11011001",  -- 7: ** **  *
    "11011111",  -- 8: ** *****
    "01101110",  -- 9:  ** *** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xBD
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01101100",  -- 4:  ** **  
    "11011010",  -- 5: ** ** * 
    "11011110",  -- 6: ** **** 
    "11011000",  -- 7: ** **   
    "11011010",  -- 8: ** ** * 
    "01101100",  -- 9:  ** **  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xBE
    "01100110",  -- 0:  **  ** 
    "01100110",  -- 1:  **  ** 
    "00000000",  -- 2:         
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "00111100",  -- 5:   ****  
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xBF
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00110000",  -- 3:   **    
    "00110000",  -- 4:   **    
    "00000000",  -- 5:         
    "00110000",  -- 6:   **    
    "00110000",  -- 7:   **    
    "01100000",  -- 8:  **     
    "11000110",  -- 9: **   ** 
    "11000110",  -- A: **   ** 
    "01111100",  -- B:  *****  
      -- Char Code: 0xC0
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111111",  -- 2: ********
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xC1
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xC2
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00011111",  -- 5:    *****
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xC3
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011111",  -- 5:    *****
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xC4
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xC5
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xC6
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00011111",  -- 5:    *****
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xC7
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "00011111",  -- 5:    *****
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xC8
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "11111000",  -- 5: *****   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xC9
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "11111000",  -- 5: *****   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xCA
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "11111111",  -- 5: ********
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xCB
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "11111111",  -- 5: ********
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xCC
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "11111000",  -- 5: *****   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xCD
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "11111000",  -- 5: *****   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xCE
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "11111111",  -- 5: ********
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xCF
    "00011000",  -- 0:    **   
    "00011000",  -- 1:    **   
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00011000",  -- 4:    **   
    "11111111",  -- 5: ********
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00011000",  -- B:    **   
      -- Char Code: 0xD0
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "11111111",  -- 7: ********
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xD1
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "01101100",  -- 4:  ** **  
    "01101100",  -- 5:  ** **  
    "01111100",  -- 6:  *****  
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xD2
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00111111",  -- 4:   ******
    "00110000",  -- 5:   **    
    "00111111",  -- 6:   ******
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xD3
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "01101111",  -- 4:  ** ****
    "01100000",  -- 5:  **     
    "01111111",  -- 6:  *******
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xD4
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "01101100",  -- 5:  ** **  
    "01101100",  -- 6:  ** **  
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xD5
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "01101100",  -- 4:  ** **  
    "01101100",  -- 5:  ** **  
    "01101100",  -- 6:  ** **  
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xD6
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111111",  -- 4:  *******
    "01100000",  -- 5:  **     
    "01101111",  -- 6:  ** ****
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xD7
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "01101111",  -- 4:  ** ****
    "01100000",  -- 5:  **     
    "01101111",  -- 6:  ** ****
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xD8
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111100",  -- 4: ******  
    "00001100",  -- 5:     **  
    "11111100",  -- 6: ******  
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xD9
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "11101100",  -- 4: *** **  
    "00001100",  -- 5:     **  
    "11111100",  -- 6: ******  
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xDA
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111111",  -- 4: ********
    "00000000",  -- 5:         
    "11111111",  -- 6: ********
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xDB
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "11101111",  -- 4: *** ****
    "00000000",  -- 5:         
    "11111111",  -- 6: ********
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xDC
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111100",  -- 4: ******  
    "00001100",  -- 5:     **  
    "11101100",  -- 6: *** **  
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xDD
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "11101100",  -- 4: *** **  
    "00001100",  -- 5:     **  
    "11101100",  -- 6: *** **  
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xDE
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111111",  -- 4: ********
    "00000000",  -- 5:         
    "11101111",  -- 6: *** ****
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xDF
    "01101100",  -- 0:  ** **  
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "01101100",  -- 3:  ** **  
    "11101111",  -- 4: *** ****
    "00000000",  -- 5:         
    "11101111",  -- 6: *** ****
    "01101100",  -- 7:  ** **  
    "01101100",  -- 8:  ** **  
    "01101100",  -- 9:  ** **  
    "01101100",  -- A:  ** **  
    "01101100",  -- B:  ** **  
      -- Char Code: 0xE0
    "01100000",  -- 0:  **     
    "00110000",  -- 1:   **    
    "00011000",  -- 2:    **   
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE1
    "00011000",  -- 0:    **   
    "00110000",  -- 1:   **    
    "01100000",  -- 2:  **     
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE2
    "00110000",  -- 0:   **    
    "01111000",  -- 1:  ****   
    "11001100",  -- 2: **  **  
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE3
    "00000000",  -- 0:         
    "01110110",  -- 1:  *** ** 
    "11011100",  -- 2: ** ***  
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE4
    "00000000",  -- 0:         
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE5
    "00111000",  -- 0:   ***   
    "01101100",  -- 1:  ** **  
    "00111000",  -- 2:   ***   
    "00000000",  -- 3:         
    "01111000",  -- 4:  ****   
    "00001100",  -- 5:     **  
    "01111100",  -- 6:  *****  
    "11001100",  -- 7: **  **  
    "11011100",  -- 8: ** ***  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE6
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01111110",  -- 3:  ****** 
    "11011011",  -- 4: ** ** **
    "00011011",  -- 5:    ** **
    "01111111",  -- 6:  *******
    "11011000",  -- 7: ** **   
    "11011011",  -- 8: ** ** **
    "01111110",  -- 9:  ****** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE7
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01111100",  -- 3:  *****  
    "11000110",  -- 4: **   ** 
    "11000000",  -- 5: **      
    "11000000",  -- 6: **      
    "11000110",  -- 7: **   ** 
    "01111100",  -- 8:  *****  
    "00011000",  -- 9:    **   
    "01101100",  -- A:  ** **  
    "00111000",  -- B:   ***   
      -- Char Code: 0xE8
    "00110000",  -- 0:   **    
    "00011000",  -- 1:    **   
    "00001100",  -- 2:     **  
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11111110",  -- 6: ******* 
    "11000000",  -- 7: **      
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xE9
    "00001100",  -- 0:     **  
    "00011000",  -- 1:    **   
    "00110000",  -- 2:   **    
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11111110",  -- 6: ******* 
    "11000000",  -- 7: **      
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xEA
    "00010000",  -- 0:    *    
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11111110",  -- 6: ******* 
    "11000000",  -- 7: **      
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xEB
    "00000000",  -- 0:         
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11111110",  -- 6: ******* 
    "11000000",  -- 7: **      
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xEC
    "01100000",  -- 0:  **     
    "00110000",  -- 1:   **    
    "00011000",  -- 2:    **   
    "00000000",  -- 3:         
    "00111000",  -- 4:   ***   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xED
    "00001100",  -- 0:     **  
    "00011000",  -- 1:    **   
    "00110000",  -- 2:   **    
    "00000000",  -- 3:         
    "00111000",  -- 4:   ***   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xEE
    "00011000",  -- 0:    **   
    "00111100",  -- 1:   ****  
    "01100110",  -- 2:  **  ** 
    "00000000",  -- 3:         
    "00111000",  -- 4:   ***   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xEF
    "00000000",  -- 0:         
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "00000000",  -- 3:         
    "00111000",  -- 4:   ***   
    "00011000",  -- 5:    **   
    "00011000",  -- 6:    **   
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00111100",  -- 9:   ****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF0
    "01111000",  -- 0:  ****   
    "00110000",  -- 1:   **    
    "01111000",  -- 2:  ****   
    "00001100",  -- 3:     **  
    "01111110",  -- 4:  ****** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF1
    "00000000",  -- 0:         
    "01110110",  -- 1:  *** ** 
    "11011100",  -- 2: ** ***  
    "00000000",  -- 3:         
    "11011100",  -- 4: ** ***  
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "01100110",  -- 7:  **  ** 
    "01100110",  -- 8:  **  ** 
    "01100110",  -- 9:  **  ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF2
    "01100000",  -- 0:  **     
    "00110000",  -- 1:   **    
    "00011000",  -- 2:    **   
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF3
    "00001100",  -- 0:     **  
    "00011000",  -- 1:    **   
    "00110000",  -- 2:   **    
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF4
    "00010000",  -- 0:    *    
    "00111000",  -- 1:   ***   
    "01101100",  -- 2:  ** **  
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF5
    "00000000",  -- 0:         
    "01110110",  -- 1:  *** ** 
    "11011100",  -- 2: ** ***  
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF6
    "00000000",  -- 0:         
    "01101100",  -- 1:  ** **  
    "01101100",  -- 2:  ** **  
    "00000000",  -- 3:         
    "01111100",  -- 4:  *****  
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11000110",  -- 7: **   ** 
    "11000110",  -- 8: **   ** 
    "01111100",  -- 9:  *****  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF7
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00011000",  -- 2:    **   
    "00011000",  -- 3:    **   
    "00000000",  -- 4:         
    "01111110",  -- 5:  ****** 
    "00000000",  -- 6:         
    "00011000",  -- 7:    **   
    "00011000",  -- 8:    **   
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF8
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "01111110",  -- 4:  ****** 
    "11001110",  -- 5: **  *** 
    "11011110",  -- 6: ** **** 
    "11110110",  -- 7: **** ** 
    "11100110",  -- 8: ***  ** 
    "11111100",  -- 9: ******  
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xF9
    "11000000",  -- 0: **      
    "01100000",  -- 1:  **     
    "00110000",  -- 2:   **    
    "00000000",  -- 3:         
    "11001100",  -- 4: **  **  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xFA
    "00001100",  -- 0:     **  
    "00011000",  -- 1:    **   
    "00110000",  -- 2:   **    
    "00000000",  -- 3:         
    "11001100",  -- 4: **  **  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xFB
    "00110000",  -- 0:   **    
    "01111000",  -- 1:  ****   
    "11001100",  -- 2: **  **  
    "00000000",  -- 3:         
    "11001100",  -- 4: **  **  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xFC
    "00000000",  -- 0:         
    "11001100",  -- 1: **  **  
    "11001100",  -- 2: **  **  
    "00000000",  -- 3:         
    "11001100",  -- 4: **  **  
    "11001100",  -- 5: **  **  
    "11001100",  -- 6: **  **  
    "11001100",  -- 7: **  **  
    "11001100",  -- 8: **  **  
    "01110110",  -- 9:  *** ** 
    "00000000",  -- A:         
    "00000000",  -- B:         
      -- Char Code: 0xFD
    "00001100",  -- 0:     **  
    "00011000",  -- 1:    **   
    "00110000",  -- 2:   **    
    "00000000",  -- 3:         
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11001110",  -- 7: **  *** 
    "01110110",  -- 8:  *** ** 
    "00000110",  -- 9:      ** 
    "11000110",  -- A: **   ** 
    "01111100",  -- B:  *****  
      -- Char Code: 0xFE
    "00000000",  -- 0:         
    "11110000",  -- 1: ****    
    "01100000",  -- 2:  **     
    "01100000",  -- 3:  **     
    "01111000",  -- 4:  ****   
    "01101100",  -- 5:  ** **  
    "01101100",  -- 6:  ** **  
    "01101100",  -- 7:  ** **  
    "01111000",  -- 8:  ****   
    "01100000",  -- 9:  **     
    "01100000",  -- A:  **     
    "11110000",  -- B: ****    
      -- Char Code: 0xFF
    "00000000",  -- 0:         
    "11000110",  -- 1: **   ** 
    "11000110",  -- 2: **   ** 
    "00000000",  -- 3:         
    "11000110",  -- 4: **   ** 
    "11000110",  -- 5: **   ** 
    "11000110",  -- 6: **   ** 
    "11001110",  -- 7: **  *** 
    "01110110",  -- 8:  *** ** 
    "00000110",  -- 9:      ** 
    "11000110",  -- A: **   ** 
    "01111100",  -- B:  *****  
    others => "00000000"
  );

  constant FONT_8X12X256 : Font_type := (
    ID       => 1,
    Width    => 8,
    Height   => 12,
    NumChars => 256,
    Data     => FONT_ROM_8X12X256
  );
  

  -- This next font table was borrowed from the Papilio Playground -- vga_text project
   constant FONT_ROM_8X16X128 : FontRom_type := (
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x01
		"00000000", -- 0
		"00000000", -- 1
		"01111110", -- 2  ******
		"10000001", -- 3 *      *
		"10100101", -- 4 * *  * *
		"10000001", -- 5 *      *
		"10000001", -- 6 *      *
		"10111101", -- 7 * **** *
		"10011001", -- 8 *  **  *
		"10000001", -- 9 *      *
		"10000001", -- a *      *
		"01111110", -- b  ******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x02
		"00000000", -- 0
		"00000000", -- 1
		"01111110", -- 2  ******
		"11111111", -- 3 ********
		"11011011", -- 4 ** ** **
		"11111111", -- 5 ********
		"11111111", -- 6 ********
		"11000011", -- 7 **    **
		"11100111", -- 8 ***  ***
		"11111111", -- 9 ********
		"11111111", -- a ********
		"01111110", -- b  ******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x03
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"01101100", -- 4  ** **
		"11111110", -- 5 *******
		"11111110", -- 6 *******
		"11111110", -- 7 *******
		"11111110", -- 8 *******
		"01111100", -- 9  *****
		"00111000", -- a   ***
		"00010000", -- b    *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x04
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00010000", -- 4    *
		"00111000", -- 5   ***
		"01111100", -- 6  *****
		"11111110", -- 7 *******
		"01111100", -- 8  *****
		"00111000", -- 9   ***
		"00010000", -- a    *
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x05
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00111100", -- 4   ****
		"00111100", -- 5   ****
		"11100111", -- 6 ***  ***
		"11100111", -- 7 ***  ***
		"11100111", -- 8 ***  ***
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x06
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00111100", -- 4   ****
		"01111110", -- 5  ******
		"11111111", -- 6 ********
		"11111111", -- 7 ********
		"01111110", -- 8  ******
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x07
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00011000", -- 6    **
		"00111100", -- 7   ****
		"00111100", -- 8   ****
		"00011000", -- 9    **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x08
		"11111111", -- 0 ********
		"11111111", -- 1 ********
		"11111111", -- 2 ********
		"11111111", -- 3 ********
		"11111111", -- 4 ********
		"11111111", -- 5 ********
		"11100111", -- 6 ***  ***
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"11100111", -- 9 ***  ***
		"11111111", -- a ********
		"11111111", -- b ********
		"11111111", -- c ********
		"11111111", -- d ********
		"11111111", -- e ********
		"11111111", -- f ********
		-- code x09
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00111100", -- 5   ****
		"01100110", -- 6  **  **
		"01000010", -- 7  *    *
		"01000010", -- 8  *    *
		"01100110", -- 9  **  **
		"00111100", -- a   ****
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0a
		"11111111", -- 0 ********
		"11111111", -- 1 ********
		"11111111", -- 2 ********
		"11111111", -- 3 ********
		"11111111", -- 4 ********
		"11000011", -- 5 **    **
		"10011001", -- 6 *  **  *
		"10111101", -- 7 * **** *
		"10111101", -- 8 * **** *
		"10011001", -- 9 *  **  *
		"11000011", -- a **    **
		"11111111", -- b ********
		"11111111", -- c ********
		"11111111", -- d ********
		"11111111", -- e ********
		"11111111", -- f ********
		-- code x0b
		"00000000", -- 0
		"00000000", -- 1
		"00011110", -- 2    ****
		"00001110", -- 3     ***
		"00011010", -- 4    ** *
		"00110010", -- 5   **  *
		"01111000", -- 6  ****
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0c
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"00111100", -- 7   ****
		"00011000", -- 8    **
		"01111110", -- 9  ******
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0d
		"00000000", -- 0
		"00000000", -- 1
		"00111111", -- 2   ******
		"00110011", -- 3   **  **
		"00111111", -- 4   ******
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"01110000", -- 9  ***
		"11110000", -- a ****
		"11100000", -- b ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0e
		"00000000", -- 0
		"00000000", -- 1
		"01111111", -- 2  *******
		"01100011", -- 3  **   **
		"01111111", -- 4  *******
		"01100011", -- 5  **   **
		"01100011", -- 6  **   **
		"01100011", -- 7  **   **
		"01100011", -- 8  **   **
		"01100111", -- 9  **  ***
		"11100111", -- a ***  ***
		"11100110", -- b ***  **
		"11000000", -- c **
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00011000", -- 4    **
		"11011011", -- 5 ** ** **
		"00111100", -- 6   ****
		"11100111", -- 7 ***  ***
		"00111100", -- 8   ****
		"11011011", -- 9 ** ** **
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x10
		"00000000", -- 0
		"10000000", -- 1 *
		"11000000", -- 2 **
		"11100000", -- 3 ***
		"11110000", -- 4 ****
		"11111000", -- 5 *****
		"11111110", -- 6 *******
		"11111000", -- 7 *****
		"11110000", -- 8 ****
		"11100000", -- 9 ***
		"11000000", -- a **
		"10000000", -- b *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x11
		"00000000", -- 0
		"00000010", -- 1       *
		"00000110", -- 2      **
		"00001110", -- 3     ***
		"00011110", -- 4    ****
		"00111110", -- 5   *****
		"11111110", -- 6 *******
		"00111110", -- 7   *****
		"00011110", -- 8    ****
		"00001110", -- 9     ***
		"00000110", -- a      **
		"00000010", -- b       *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x12
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"01111110", -- 4  ******
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"01111110", -- 8  ******
		"00111100", -- 9   ****
		"00011000", -- a    **
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x13
		"00000000", -- 0
		"00000000", -- 1
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"00000000", -- 9
		"01100110", -- a  **  **
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x14
		"00000000", -- 0
		"00000000", -- 1
		"01111111", -- 2  *******
		"11011011", -- 3 ** ** **
		"11011011", -- 4 ** ** **
		"11011011", -- 5 ** ** **
		"01111011", -- 6  **** **
		"00011011", -- 7    ** **
		"00011011", -- 8    ** **
		"00011011", -- 9    ** **
		"00011011", -- a    ** **
		"00011011", -- b    ** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x15
		"00000000", -- 0
		"01111100", -- 1  *****
		"11000110", -- 2 **   **
		"01100000", -- 3  **
		"00111000", -- 4   ***
		"01101100", -- 5  ** **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"01101100", -- 8  ** **
		"00111000", -- 9   ***
		"00001100", -- a     **
		"11000110", -- b **   **
		"01111100", -- c  *****
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x16
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"11111110", -- 8 *******
		"11111110", -- 9 *******
		"11111110", -- a *******
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x17
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"01111110", -- 4  ******
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"01111110", -- 8  ******
		"00111100", -- 9   ****
		"00011000", -- a    **
		"01111110", -- b  ******
		"00110000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x18
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"01111110", -- 4  ******
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x19
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"01111110", -- 9  ******
		"00111100", -- a   ****
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00011000", -- 5    **
		"00001100", -- 6     **
		"11111110", -- 7 *******
		"00001100", -- 8     **
		"00011000", -- 9    **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00110000", -- 5   **
		"01100000", -- 6  **
		"11111110", -- 7 *******
		"01100000", -- 8  **
		"00110000", -- 9   **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"11000000", -- 6 **
		"11000000", -- 7 **
		"11000000", -- 8 **
		"11111110", -- 9 *******
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00100100", -- 5   *  *
		"01100110", -- 6  **  **
		"11111111", -- 7 ********
		"01100110", -- 8  **  **
		"00100100", -- 9   *  *
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00010000", -- 4    *
		"00111000", -- 5   ***
		"00111000", -- 6   ***
		"01111100", -- 7  *****
		"01111100", -- 8  *****
		"11111110", -- 9 *******
		"11111110", -- a *******
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"11111110", -- 4 *******
		"11111110", -- 5 *******
		"01111100", -- 6  *****
		"01111100", -- 7  *****
		"00111000", -- 8   ***
		"00111000", -- 9   ***
		"00010000", -- a    *
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x20
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x21
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"00111100", -- 4   ****
		"00111100", -- 5   ****
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00000000", -- 9
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x22
		"00000000", -- 0
		"01100110", -- 1  **  **
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"00100100", -- 4   *  *
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x23
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"01101100", -- 3  ** **
		"01101100", -- 4  ** **
		"11111110", -- 5 *******
		"01101100", -- 6  ** **
		"01101100", -- 7  ** **
		"01101100", -- 8  ** **
		"11111110", -- 9 *******
		"01101100", -- a  ** **
		"01101100", -- b  ** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x24
		"00011000", -- 0     **
		"00011000", -- 1     **
		"01111100", -- 2   *****
		"11000110", -- 3  **   **
		"11000010", -- 4  **    *
		"11000000", -- 5  **
		"01111100", -- 6   *****
		"00000110", -- 7       **
		"00000110", -- 8       **
		"10000110", -- 9  *    **
		"11000110", -- a  **   **
		"01111100", -- b   *****
		"00011000", -- c     **
		"00011000", -- d     **
		"00000000", -- e
		"00000000", -- f
		-- code x25
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"11000010", -- 4 **    *
		"11000110", -- 5 **   **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"01100000", -- 9  **
		"11000110", -- a **   **
		"10000110", -- b *    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x26
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01101100", -- 3  ** **
		"01101100", -- 4  ** **
		"00111000", -- 5   ***
		"01110110", -- 6  *** **
		"11011100", -- 7 ** ***
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x27
		"00000000", -- 0
		"00110000", -- 1   **
		"00110000", -- 2   **
		"00110000", -- 3   **
		"01100000", -- 4  **
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x28
		"00000000", -- 0
		"00000000", -- 1
		"00001100", -- 2     **
		"00011000", -- 3    **
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00011000", -- a    **
		"00001100", -- b     **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x29
		"00000000", -- 0
		"00000000", -- 1
		"00110000", -- 2   **
		"00011000", -- 3    **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00001100", -- 7     **
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00011000", -- a    **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01100110", -- 5  **  **
		"00111100", -- 6   ****
		"11111111", -- 7 ********
		"00111100", -- 8   ****
		"01100110", -- 9  **  **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00011000", -- 5    **
		"00011000", -- 6    **
		"01111110", -- 7  ******
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00011000", -- 9    **
		"00011000", -- a    **
		"00011000", -- b    **
		"00110000", -- c   **
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"01111110", -- 7  ******
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000010", -- 4       *
		"00000110", -- 5      **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"01100000", -- 9  **
		"11000000", -- a **
		"10000000", -- b *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x30
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11001110", -- 5 **  ***
		"11011110", -- 6 ** ****
		"11110110", -- 7 **** **
		"11100110", -- 8 ***  **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x31
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2
		"00111000", -- 3
		"01111000", -- 4    **
		"00011000", -- 5   ***
		"00011000", -- 6  ****
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"01111110", -- b    **
		"00000000", -- c    **
		"00000000", -- d  ******
		"00000000", -- e
		"00000000", -- f
		-- code x32
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		"01100000", -- 8  **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x33
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00000110", -- 5      **
		"00111100", -- 6   ****
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x34
		"00000000", -- 0
		"00000000", -- 1
		"00001100", -- 2     **
		"00011100", -- 3    ***
		"00111100", -- 4   ****
		"01101100", -- 5  ** **
		"11001100", -- 6 **  **
		"11111110", -- 7 *******
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00001100", -- a     **
		"00011110", -- b    ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x35
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"11000000", -- 3 **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11111100", -- 6 ******
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x36
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01100000", -- 3  **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11111100", -- 6 ******
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x37
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00000110", -- 5      **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110000", -- a   **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x38
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"01111100", -- 6  *****
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x39
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"01111110", -- 6  ******
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"00001100", -- a     **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00011000", -- 9    **
		"00011000", -- a    **
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00011000", -- 9    **
		"00011000", -- a    **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000110", -- 3      **
		"00001100", -- 4     **
		"00011000", -- 5    **
		"00110000", -- 6   **
		"01100000", -- 7  **
		"00110000", -- 8   **
		"00011000", -- 9    **
		"00001100", -- a     **
		"00000110", -- b      **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111110", -- 5  ******
		"00000000", -- 6
		"00000000", -- 7
		"01111110", -- 8  ******
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"01100000", -- 3  **
		"00110000", -- 4   **
		"00011000", -- 5    **
		"00001100", -- 6     **
		"00000110", -- 7      **
		"00001100", -- 8     **
		"00011000", -- 9    **
		"00110000", -- a   **
		"01100000", -- b  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3f
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00000000", -- 9
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x40
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11011110", -- 6 ** ****
		"11011110", -- 7 ** ****
		"11011110", -- 8 ** ****
		"11011100", -- 9 ** ***
		"11000000", -- a **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x41
		"00000000", -- 0
		"00000000", -- 1
		"00010000", -- 2    *
		"00111000", -- 3   ***
		"01101100", -- 4  ** **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11111110", -- 7 *******
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"11000110", -- b **   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x42
		"00000000", -- 0
		"00000000", -- 1
		"11111100", -- 2 ******
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01111100", -- 6  *****
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11111100", -- b ******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x43
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"11000010", -- 4 **    *
		"11000000", -- 5 **
		"11000000", -- 6 **
		"11000000", -- 7 **
		"11000000", -- 8 **
		"11000010", -- 9 **    *
		"01100110", -- a  **  **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x44
		"00000000", -- 0
		"00000000", -- 1
		"11111000", -- 2 *****
		"01101100", -- 3  ** **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01101100", -- a  ** **
		"11111000", -- b *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x45
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"01100110", -- 3  **  **
		"01100010", -- 4  **   *
		"01101000", -- 5  ** *
		"01111000", -- 6  ****
		"01101000", -- 7  ** *
		"01100000", -- 8  **
		"01100010", -- 9  **   *
		"01100110", -- a  **  **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x46
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"01100110", -- 3  **  **
		"01100010", -- 4  **   *
		"01101000", -- 5  ** *
		"01111000", -- 6  ****
		"01101000", -- 7  ** *
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x47
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"11000010", -- 4 **    *
		"11000000", -- 5 **
		"11000000", -- 6 **
		"11011110", -- 7 ** ****
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"01100110", -- a  **  **
		"00111010", -- b   *** *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x48
		"00000000", -- 0
		"00000000", -- 1
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11111110", -- 6 *******
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"11000110", -- b **   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x49
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x4a
		"00000000", -- 0
		"00000000", -- 1
		"00011110", -- 2    ****
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00001100", -- 7     **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x4b
		"00000000", -- 0
		"00000000", -- 1
		"11100110", -- 2 ***  **
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01101100", -- 5  ** **
		"01111000", -- 6  ****
		"01111000", -- 7  ****
		"01101100", -- 8  ** **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x4c
		"00000000", -- 0
		"00000000", -- 1
		"11110000", -- 2 ****
		"01100000", -- 3  **
		"01100000", -- 4  **
		"01100000", -- 5  **
		"01100000", -- 6  **
		"01100000", -- 7  **
		"01100000", -- 8  **
		"01100010", -- 9  **   *
		"01100110", -- a  **  **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x4d
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11100111", -- 3 ***  ***
		"11111111", -- 4 ********
		"11111111", -- 5 ********
		"11011011", -- 6 ** ** **
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"11000011", -- 9 **    **
		"11000011", -- a **    **
		"11000011", -- b **    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x4e
		"00000000", -- 0
		"00000000", -- 1
		"11000110", -- 2 **   **
		"11100110", -- 3 ***  **
		"11110110", -- 4 **** **
		"11111110", -- 5 *******
		"11011110", -- 6 ** ****
		"11001110", -- 7 **  ***
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"11000110", -- b **   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x4f
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x50
		"00000000", -- 0
		"00000000", -- 1
		"11111100", -- 2 ******
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01111100", -- 6  *****
		"01100000", -- 7  **
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x510
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11010110", -- 9 ** * **
		"11011110", -- a ** ****
		"01111100", -- b  *****
		"00001100", -- c     **
		"00001110", -- d     ***
		"00000000", -- e
		"00000000", -- f
		-- code x52
		"00000000", -- 0
		"00000000", -- 1
		"11111100", -- 2 ******
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01111100", -- 6  *****
		"01101100", -- 7  ** **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x53
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"01100000", -- 5  **
		"00111000", -- 6   ***
		"00001100", -- 7     **
		"00000110", -- 8      **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x54
		"00000000", -- 0
		"00000000", -- 1
		"11111111", -- 2 ********
		"11011011", -- 3 ** ** **
		"10011001", -- 4 *  **  *
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x55
		"00000000", -- 0
		"00000000", -- 1
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x56
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"01100110", -- 9  **  **
		"00111100", -- a   ****
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x57
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11011011", -- 7 ** ** **
		"11011011", -- 8 ** ** **
		"11111111", -- 9 ********
		"01100110", -- a  **  **
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f

		-- code x58
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"01100110", -- 4  **  **
		"00111100", -- 5   ****
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00111100", -- 8   ****
		"01100110", -- 9  **  **
		"11000011", -- a **    **
		"11000011", -- b **    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x59
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"01100110", -- 5  **  **
		"00111100", -- 6   ****
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5a
		"00000000", -- 0
		"00000000", -- 1
		"11111111", -- 2 ********
		"11000011", -- 3 **    **
		"10000110", -- 4 *    **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		"01100000", -- 8  **
		"11000001", -- 9 **     *
		"11000011", -- a **    **
		"11111111", -- b ********
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5b
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"00110000", -- 3   **
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110000", -- a   **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"10000000", -- 3 *
		"11000000", -- 4 **
		"11100000", -- 5 ***
		"01110000", -- 6  ***
		"00111000", -- 7   ***
		"00011100", -- 8    ***
		"00001110", -- 9     ***
		"00000110", -- a      **
		"00000010", -- b       *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5d
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00001100", -- 7     **
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00001100", -- a     **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5e
		"00010000", -- 0    *
		"00111000", -- 1   ***
		"01101100", -- 2  ** **
		"11000110", -- 3 **   **
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"11111111", -- d ********
		"00000000", -- e
		"00000000", -- f
		-- code x60
		"00110000", -- 0   **
		"00110000", -- 1   **
		"00011000", -- 2    **
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x61
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111000", -- 5  ****
		"00001100", -- 6     **
		"01111100", -- 7  *****
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x62
		"00000000", -- 0
		"00000000", -- 1
		"11100000", -- 2  ***
		"01100000", -- 3   **
		"01100000", -- 4   **
		"01111000", -- 5   ****
		"01101100", -- 6   ** **
		"01100110", -- 7   **  **
		"01100110", -- 8   **  **
		"01100110", -- 9   **  **
		"01100110", -- a   **  **
		"01111100", -- b   *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x63
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"11000000", -- 7 **
		"11000000", -- 8 **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x64
		"00000000", -- 0
		"00000000", -- 1
		"00011100", -- 2    ***
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00111100", -- 5   ****
		"01101100", -- 6  ** **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x65
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"11111110", -- 7 *******
		"11000000", -- 8 **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x66
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01101100", -- 3  ** **
		"01100100", -- 4  **  *
		"01100000", -- 5  **
		"11110000", -- 6 ****
		"01100000", -- 7  **
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x67
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01110110", -- 5  *** **
		"11001100", -- 6 **  **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111100", -- b  *****
		"00001100", -- c     **
		"11001100", -- d **  **
		"01111000", -- e  ****
		"00000000", -- f
		-- code x68
		"00000000", -- 0
		"00000000", -- 1
		"11100000", -- 2 ***
		"01100000", -- 3  **
		"01100000", -- 4  **
		"01101100", -- 5  ** **
		"01110110", -- 6  *** **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x69
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00000000", -- 4
		"00111000", -- 5   ***
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x6a
		"00000000", -- 0
		"00000000", -- 1
		"00000110", -- 2      **
		"00000110", -- 3      **
		"00000000", -- 4
		"00001110", -- 5     ***
		"00000110", -- 6      **
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"00000110", -- a      **
		"00000110", -- b      **
		"01100110", -- c  **  **
		"01100110", -- d  **  **
		"00111100", -- e   ****
		"00000000", -- f
		-- code x6b
		"00000000", -- 0
		"00000000", -- 1
		"11100000", -- 2 ***
		"01100000", -- 3  **
		"01100000", -- 4  **
		"01100110", -- 5  **  **
		"01101100", -- 6  ** **
		"01111000", -- 7  ****
		"01111000", -- 8  ****
		"01101100", -- 9  ** **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x6c
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x6d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11100110", -- 5 ***  **
		"11111111", -- 6 ********
		"11011011", -- 7 ** ** **
		"11011011", -- 8 ** ** **
		"11011011", -- 9 ** ** **
		"11011011", -- a ** ** **
		"11011011", -- b ** ** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x6e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11011100", -- 5 ** ***
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x6f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x70
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11011100", -- 5 ** ***
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"01111100", -- b  *****
		"01100000", -- c  **
		"01100000", -- d  **
		"11110000", -- e ****
		"00000000", -- f
		-- code x71
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01110110", -- 5  *** **
		"11001100", -- 6 **  **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111100", -- b  *****
		"00001100", -- c     **
		"00001100", -- d     **
		"00011110", -- e    ****
		"00000000", -- f
		-- code x72
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11011100", -- 5 ** ***
		"01110110", -- 6  *** **
		"01100110", -- 7  **  **
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x73
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"01100000", -- 7  **
		"00111000", -- 8   ***
		"00001100", -- 9     **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x74
		"00000000", -- 0
		"00000000", -- 1
		"00010000", -- 2    *
		"00110000", -- 3   **
		"00110000", -- 4   **
		"11111100", -- 5 ******
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110110", -- a   ** **
		"00011100", -- b    ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x75
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11001100", -- 5 **  **
		"11001100", -- 6 **  **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x76
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"01100110", -- 9  **  **
		"00111100", -- a   ****
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x77
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11000011", -- 7 **    **
		"11011011", -- 8 ** ** **
		"11011011", -- 9 ** ** **
		"11111111", -- a ********
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x78
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000011", -- 5 **    **
		"01100110", -- 6  **  **
		"00111100", -- 7   ****
		"00011000", -- 8    **
		"00111100", -- 9   ****
		"01100110", -- a  **  **
		"11000011", -- b **    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x79
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111110", -- b  ******
		"00000110", -- c      **
		"00001100", -- d     **
		"11111000", -- e *****
		"00000000", -- f
		-- code x7a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11111110", -- 5 *******
		"11001100", -- 6 **  **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"01100000", -- 9  **
		"11000110", -- a **   **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7b
		"00000000", -- 0
		"00000000", -- 1
		"00001110", -- 2     ***
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"01110000", -- 6  ***
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00001110", -- b     ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7c
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00000000", -- 6
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7d
		"00000000", -- 0
		"00000000", -- 1
		"01110000", -- 2  ***
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00001110", -- 6     ***
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"01110000", -- b  ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7e
		"00000000", -- 0
		"00000000", -- 1
		"01110110", -- 2  *** **
		"11011100", -- 3 ** ***
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00010000", -- 4    *
		"00111000", -- 5   ***
		"01101100", -- 6  ** **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11111110", -- a *******
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
    others => "00000000"
  );

  constant FONT_8X16X128 : Font_type := (
    ID       => 2,
    Width    => 8,
    Height   => 16,
    NumChars => 128,
    Data     => FONT_ROM_8X16X128
  );
  
 constant FONT_ROM_8X16X128_2 : FontRom_type := (
       -- Char Code: 0x00
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x01
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "11111111",  -- 3: ********
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "11111111",  -- 6: ********
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "11111111",  -- 9: ********
    "00000000",  -- A:         
    "00000000",  -- B:         
    "11111111",  -- C: ********
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x02
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111111",  -- 2: ********
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "11111111",  -- 5: ********
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "11111111",  -- 8: ********
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "11111111",  -- B: ********
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x03
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00100100",  -- 2:   *  *  
    "00100100",  -- 3:   *  *  
    "00100100",  -- 4:   *  *  
    "00100100",  -- 5:   *  *  
    "00100100",  -- 6:   *  *  
    "00100100",  -- 7:   *  *  
    "00100100",  -- 8:   *  *  
    "00100100",  -- 9:   *  *  
    "00100100",  -- A:   *  *  
    "00100100",  -- B:   *  *  
    "00100100",  -- C:   *  *  
    "00100100",  -- D:   *  *  
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x04
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01001001",  -- 2:  *  *  *
    "01001001",  -- 3:  *  *  *
    "01001001",  -- 4:  *  *  *
    "01001001",  -- 5:  *  *  *
    "01001001",  -- 6:  *  *  *
    "01001001",  -- 7:  *  *  *
    "01001001",  -- 8:  *  *  *
    "01001001",  -- 9:  *  *  *
    "01001001",  -- A:  *  *  *
    "01001001",  -- B:  *  *  *
    "01001001",  -- C:  *  *  *
    "01001001",  -- D:  *  *  *
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x05
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10010010",  -- 2: *  *  * 
    "10010010",  -- 3: *  *  * 
    "10010010",  -- 4: *  *  * 
    "10010010",  -- 5: *  *  * 
    "10010010",  -- 6: *  *  * 
    "10010010",  -- 7: *  *  * 
    "10010010",  -- 8: *  *  * 
    "10010010",  -- 9: *  *  * 
    "10010010",  -- A: *  *  * 
    "10010010",  -- B: *  *  * 
    "10010010",  -- C: *  *  * 
    "10010010",  -- D: *  *  * 
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x06
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01010101",  -- 2:  * * * *
    "01010101",  -- 3:  * * * *
    "01010101",  -- 4:  * * * *
    "01010101",  -- 5:  * * * *
    "01010101",  -- 6:  * * * *
    "01010101",  -- 7:  * * * *
    "01010101",  -- 8:  * * * *
    "01010101",  -- 9:  * * * *
    "01010101",  -- A:  * * * *
    "01010101",  -- B:  * * * *
    "01010101",  -- C:  * * * *
    "01010101",  -- D:  * * * *
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x07
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10101010",  -- 2: * * * * 
    "10101010",  -- 3: * * * * 
    "10101010",  -- 4: * * * * 
    "10101010",  -- 5: * * * * 
    "10101010",  -- 6: * * * * 
    "10101010",  -- 7: * * * * 
    "10101010",  -- 8: * * * * 
    "10101010",  -- 9: * * * * 
    "10101010",  -- A: * * * * 
    "10101010",  -- B: * * * * 
    "10101010",  -- C: * * * * 
    "10101010",  -- D: * * * * 
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x08
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "11111111",  -- 3: ********
    "00000000",  -- 4:         
    "11111111",  -- 5: ********
    "00000000",  -- 6:         
    "11111111",  -- 7: ********
    "00000000",  -- 8:         
    "11111111",  -- 9: ********
    "00000000",  -- A:         
    "11111111",  -- B: ********
    "00000000",  -- C:         
    "11111111",  -- D: ********
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x09
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111100",  -- 2: ******  
    "11110011",  -- 3: ****  **
    "11111100",  -- 4: ******  
    "11110011",  -- 5: ****  **
    "11111100",  -- 6: ******  
    "11110011",  -- 7: ****  **
    "11111100",  -- 8: ******  
    "11110011",  -- 9: ****  **
    "11111100",  -- A: ******  
    "11110011",  -- B: ****  **
    "11111100",  -- C: ******  
    "11110011",  -- D: ****  **
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x0A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111111",  -- 2:   ******
    "11001111",  -- 3: **  ****
    "00111111",  -- 4:   ******
    "11001111",  -- 5: **  ****
    "00111111",  -- 6:   ******
    "11001111",  -- 7: **  ****
    "00111111",  -- 8:   ******
    "11001111",  -- 9: **  ****
    "00111111",  -- A:   ******
    "11001111",  -- B: **  ****
    "00111111",  -- C:   ******
    "11001111",  -- D: **  ****
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x0B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000011",  -- 2:       **
    "00001100",  -- 3:     **  
    "00000011",  -- 4:       **
    "00001100",  -- 5:     **  
    "00000011",  -- 6:       **
    "00001100",  -- 7:     **  
    "00000011",  -- 8:       **
    "00001100",  -- 9:     **  
    "00000011",  -- A:       **
    "00001100",  -- B:     **  
    "00000011",  -- C:       **
    "00001100",  -- D:     **  
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x0C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11000000",  -- 2: **      
    "00110000",  -- 3:   **    
    "11000000",  -- 4: **      
    "00110000",  -- 5:   **    
    "11000000",  -- 6: **      
    "00110000",  -- 7:   **    
    "11000000",  -- 8: **      
    "00110000",  -- 9:   **    
    "11000000",  -- A: **      
    "00110000",  -- B:   **    
    "11000000",  -- C: **      
    "00110000",  -- D:   **    
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x0D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01100110",  -- 3:  **  ** 
    "01100110",  -- 4:  **  ** 
    "01100110",  -- 5:  **  ** 
    "01100110",  -- 6:  **  ** 
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "01100110",  -- 9:  **  ** 
    "01100110",  -- A:  **  ** 
    "01100110",  -- B:  **  ** 
    "01100110",  -- C:  **  ** 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x0E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111111",  -- 2: ********
    "10011001",  -- 3: *  **  *
    "10011001",  -- 4: *  **  *
    "10011001",  -- 5: *  **  *
    "10011001",  -- 6: *  **  *
    "11111111",  -- 7: ********
    "11111111",  -- 8: ********
    "10011001",  -- 9: *  **  *
    "10011001",  -- A: *  **  *
    "10011001",  -- B: *  **  *
    "10011001",  -- C: *  **  *
    "11111111",  -- D: ********
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x0F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00001111",  -- 2:     ****
    "00001111",  -- 3:     ****
    "00001111",  -- 4:     ****
    "00001111",  -- 5:     ****
    "00001111",  -- 6:     ****
    "00001111",  -- 7:     ****
    "00001111",  -- 8:     ****
    "00001111",  -- 9:     ****
    "00001111",  -- A:     ****
    "00001111",  -- B:     ****
    "00001111",  -- C:     ****
    "00001111",  -- D:     ****
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x10
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11110000",  -- 2: ****    
    "11110000",  -- 3: ****    
    "11110000",  -- 4: ****    
    "11110000",  -- 5: ****    
    "11110000",  -- 6: ****    
    "11110000",  -- 7: ****    
    "11110000",  -- 8: ****    
    "11110000",  -- 9: ****    
    "11110000",  -- A: ****    
    "11110000",  -- B: ****    
    "11110000",  -- C: ****    
    "11110000",  -- D: ****    
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x11
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111111",  -- 2: ********
    "11111111",  -- 3: ********
    "11111111",  -- 4: ********
    "11111111",  -- 5: ********
    "11111111",  -- 6: ********
    "11111111",  -- 7: ********
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x12
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "11111111",  -- 8: ********
    "11111111",  -- 9: ********
    "11111111",  -- A: ********
    "11111111",  -- B: ********
    "11111111",  -- C: ********
    "11111111",  -- D: ********
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x13
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00001111",  -- 2:     ****
    "00001111",  -- 3:     ****
    "00001111",  -- 4:     ****
    "00001111",  -- 5:     ****
    "00001111",  -- 6:     ****
    "00001111",  -- 7:     ****
    "00001111",  -- 8:     ****
    "00001111",  -- 9:     ****
    "00001111",  -- A:     ****
    "00001111",  -- B:     ****
    "00001111",  -- C:     ****
    "00001111",  -- D:     ****
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x14
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11110000",  -- 2: ****    
    "11110000",  -- 3: ****    
    "11110000",  -- 4: ****    
    "11110000",  -- 5: ****    
    "11110000",  -- 6: ****    
    "11110000",  -- 7: ****    
    "11110000",  -- 8: ****    
    "11110000",  -- 9: ****    
    "11110000",  -- A: ****    
    "11110000",  -- B: ****    
    "11110000",  -- C: ****    
    "11110000",  -- D: ****    
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x15
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "01111110",  -- 3:  ****** 
    "01000010",  -- 4:  *    * 
    "01000010",  -- 5:  *    * 
    "01000010",  -- 6:  *    * 
    "01000010",  -- 7:  *    * 
    "01000010",  -- 8:  *    * 
    "01000010",  -- 9:  *    * 
    "01000010",  -- A:  *    * 
    "01000010",  -- B:  *    * 
    "01111110",  -- C:  ****** 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x16
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111111",  -- 2: ********
    "10000001",  -- 3: *      *
    "10000001",  -- 4: *      *
    "10000001",  -- 5: *      *
    "10000001",  -- 6: *      *
    "10000001",  -- 7: *      *
    "10000001",  -- 8: *      *
    "10000001",  -- 9: *      *
    "10000001",  -- A: *      *
    "10000001",  -- B: *      *
    "10000001",  -- C: *      *
    "11111111",  -- D: ********
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x17
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01001001",  -- 2:  *  *  *
    "00100100",  -- 3:   *  *  
    "01001001",  -- 4:  *  *  *
    "00100100",  -- 5:   *  *  
    "01001001",  -- 6:  *  *  *
    "00100100",  -- 7:   *  *  
    "01001001",  -- 8:  *  *  *
    "00100100",  -- 9:   *  *  
    "01001001",  -- A:  *  *  *
    "00100100",  -- B:   *  *  
    "01001001",  -- C:  *  *  *
    "00100100",  -- D:   *  *  
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x18
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10010010",  -- 2: *  *  * 
    "00100100",  -- 3:   *  *  
    "10010010",  -- 4: *  *  * 
    "00100100",  -- 5:   *  *  
    "10010010",  -- 6: *  *  * 
    "00100100",  -- 7:   *  *  
    "10010010",  -- 8: *  *  * 
    "00100100",  -- 9:   *  *  
    "10010010",  -- A: *  *  * 
    "00100100",  -- B:   *  *  
    "10010010",  -- C: *  *  * 
    "00100100",  -- D:   *  *  
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x19
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10010010",  -- 2: *  *  * 
    "01001001",  -- 3:  *  *  *
    "10010010",  -- 4: *  *  * 
    "01001001",  -- 5:  *  *  *
    "10010010",  -- 6: *  *  * 
    "01001001",  -- 7:  *  *  *
    "10010010",  -- 8: *  *  * 
    "01001001",  -- 9:  *  *  *
    "10010010",  -- A: *  *  * 
    "01001001",  -- B:  *  *  *
    "10010010",  -- C: *  *  * 
    "01001001",  -- D:  *  *  *
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x1A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10101010",  -- 2: * * * * 
    "01010101",  -- 3:  * * * *
    "10101010",  -- 4: * * * * 
    "01010101",  -- 5:  * * * *
    "10101010",  -- 6: * * * * 
    "01010101",  -- 7:  * * * *
    "10101010",  -- 8: * * * * 
    "01010101",  -- 9:  * * * *
    "10101010",  -- A: * * * * 
    "01010101",  -- B:  * * * *
    "10101010",  -- C: * * * * 
    "01010101",  -- D:  * * * *
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x1B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01010101",  -- 2:  * * * *
    "10101010",  -- 3: * * * * 
    "01010101",  -- 4:  * * * *
    "10101010",  -- 5: * * * * 
    "01010101",  -- 6:  * * * *
    "10101010",  -- 7: * * * * 
    "01010101",  -- 8:  * * * *
    "10101010",  -- 9: * * * * 
    "01010101",  -- A:  * * * *
    "10101010",  -- B: * * * * 
    "01010101",  -- C:  * * * *
    "10101010",  -- D: * * * * 
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x1C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10110110",  -- 2: * ** ** 
    "11011011",  -- 3: ** ** **
    "10110110",  -- 4: * ** ** 
    "11011011",  -- 5: ** ** **
    "10110110",  -- 6: * ** ** 
    "11011011",  -- 7: ** ** **
    "10110110",  -- 8: * ** ** 
    "11011011",  -- 9: ** ** **
    "10110110",  -- A: * ** ** 
    "11011011",  -- B: ** ** **
    "10110110",  -- C: * ** ** 
    "11011011",  -- D: ** ** **
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x1D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01101101",  -- 2:  ** ** *
    "11011011",  -- 3: ** ** **
    "01101101",  -- 4:  ** ** *
    "11011011",  -- 5: ** ** **
    "01101101",  -- 6:  ** ** *
    "11011011",  -- 7: ** ** **
    "01101101",  -- 8:  ** ** *
    "11011011",  -- 9: ** ** **
    "01101101",  -- A:  ** ** *
    "11011011",  -- B: ** ** **
    "01101101",  -- C:  ** ** *
    "11011011",  -- D: ** ** **
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x1E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01101101",  -- 2:  ** ** *
    "10110110",  -- 3: * ** ** 
    "01101101",  -- 4:  ** ** *
    "10110110",  -- 5: * ** ** 
    "01101101",  -- 6:  ** ** *
    "10110110",  -- 7: * ** ** 
    "01101101",  -- 8:  ** ** *
    "10110110",  -- 9: * ** ** 
    "01101101",  -- A:  ** ** *
    "10110110",  -- B: * ** ** 
    "01101101",  -- C:  ** ** *
    "10110110",  -- D: * ** ** 
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x1F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111111",  -- 2: ********
    "11111111",  -- 3: ********
    "11111111",  -- 4: ********
    "11111111",  -- 5: ********
    "11111111",  -- 6: ********
    "11111111",  -- 7: ********
    "11111111",  -- 8: ********
    "11111111",  -- 9: ********
    "11111111",  -- A: ********
    "11111111",  -- B: ********
    "11111111",  -- C: ********
    "11111111",  -- D: ********
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x20
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x21
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00010000",  -- 3:    *    
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x22
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01000100",  -- 2:  *   *  
    "01000100",  -- 3:  *   *  
    "01000100",  -- 4:  *   *  
    "01000100",  -- 5:  *   *  
    "01000100",  -- 6:  *   *  
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x23
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01000100",  -- 2:  *   *  
    "01000100",  -- 3:  *   *  
    "11111110",  -- 4: ******* 
    "01000100",  -- 5:  *   *  
    "01000100",  -- 6:  *   *  
    "01000100",  -- 7:  *   *  
    "01000100",  -- 8:  *   *  
    "01000100",  -- 9:  *   *  
    "11111110",  -- A: ******* 
    "01000100",  -- B:  *   *  
    "01000100",  -- C:  *   *  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x24
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10010010",  -- 3: *  *  * 
    "10010000",  -- 4: *  *    
    "10010000",  -- 5: *  *    
    "10010000",  -- 6: *  *    
    "01111100",  -- 7:  *****  
    "00010010",  -- 8:    *  * 
    "00010010",  -- 9:    *  * 
    "00010010",  -- A:    *  * 
    "10010010",  -- B: *  *  * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x25
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01100000",  -- 2:  **     
    "10010000",  -- 3: *  *    
    "10010010",  -- 4: *  *  * 
    "01100100",  -- 5:  **  *  
    "00001000",  -- 6:     *   
    "00010000",  -- 7:    *    
    "00100000",  -- 8:   *     
    "01001100",  -- 9:  *  **  
    "10010010",  -- A: *  *  * 
    "00010010",  -- B:    *  * 
    "00001100",  -- C:     **  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x26
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00110000",  -- 2:   **    
    "01001000",  -- 3:  *  *   
    "10001000",  -- 4: *   *   
    "10001000",  -- 5: *   *   
    "10010000",  -- 6: *  *    
    "01110000",  -- 7:  ***    
    "01010000",  -- 8:  * *    
    "10001010",  -- 9: *   * * 
    "10000100",  -- A: *    *  
    "10000100",  -- B: *    *  
    "01111010",  -- C:  **** * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x27
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00010000",  -- 3:    *    
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x28
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00100000",  -- 3:   *     
    "00100000",  -- 4:   *     
    "01000000",  -- 5:  *      
    "01000000",  -- 6:  *      
    "01000000",  -- 7:  *      
    "01000000",  -- 8:  *      
    "01000000",  -- 9:  *      
    "00100000",  -- A:   *     
    "00100000",  -- B:   *     
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x29
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00001000",  -- 3:     *   
    "00001000",  -- 4:     *   
    "00000100",  -- 5:      *  
    "00000100",  -- 6:      *  
    "00000100",  -- 7:      *  
    "00000100",  -- 8:      *  
    "00000100",  -- 9:      *  
    "00001000",  -- A:     *   
    "00001000",  -- B:     *   
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x2A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10010010",  -- 2: *  *  * 
    "10010010",  -- 3: *  *  * 
    "01010100",  -- 4:  * * *  
    "01010100",  -- 5:  * * *  
    "00111000",  -- 6:   ***   
    "11111110",  -- 7: ******* 
    "00111000",  -- 8:   ***   
    "01010100",  -- 9:  * * *  
    "01010100",  -- A:  * * *  
    "10010010",  -- B: *  *  * 
    "10010010",  -- C: *  *  * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x2B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00010000",  -- 3:    *    
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "11111110",  -- 7: ******* 
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x2C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00010000",  -- B:    *    
    "00100000",  -- C:   *     
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x2D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "11111110",  -- 7: ******* 
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x2E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x2F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000010",  -- 4:       * 
    "00000100",  -- 5:      *  
    "00001000",  -- 6:     *   
    "00010000",  -- 7:    *    
    "00100000",  -- 8:   *     
    "01000000",  -- 9:  *      
    "10000000",  -- A: *       
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x30
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111000",  -- 2:   ***   
    "01000100",  -- 3:  *   *  
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10001010",  -- 6: *   * * 
    "10010010",  -- 7: *  *  * 
    "10100010",  -- 8: * *   * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "01000100",  -- B:  *   *  
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x31
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00110000",  -- 3:   **    
    "01010000",  -- 4:  * *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x32
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "00000010",  -- 4:       * 
    "00000010",  -- 5:       * 
    "00000010",  -- 6:       * 
    "01111100",  -- 7:  *****  
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "11111110",  -- C: ******* 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x33
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "00000010",  -- 4:       * 
    "00000010",  -- 5:       * 
    "00000010",  -- 6:       * 
    "01111100",  -- 7:  *****  
    "00000010",  -- 8:       * 
    "00000010",  -- 9:       * 
    "00000010",  -- A:       * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x34
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00001000",  -- 2:     *   
    "00011000",  -- 3:    **   
    "00101000",  -- 4:   * *   
    "01001000",  -- 5:  *  *   
    "10001000",  -- 6: *   *   
    "10001000",  -- 7: *   *   
    "11111110",  -- 8: ******* 
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00001000",  -- B:     *   
    "00011100",  -- C:    ***  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x35
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111110",  -- 2: ******* 
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "01111100",  -- 7:  *****  
    "00000010",  -- 8:       * 
    "00000010",  -- 9:       * 
    "00000010",  -- A:       * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x36
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111110",  -- 2:  ****** 
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "01111100",  -- 7:  *****  
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x37
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111110",  -- 2: ******* 
    "00000010",  -- 3:       * 
    "00000010",  -- 4:       * 
    "00000100",  -- 5:      *  
    "00001000",  -- 6:     *   
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x38
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "01111100",  -- 7:  *****  
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x39
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "01111100",  -- 7:  *****  
    "00000010",  -- 8:       * 
    "00000010",  -- 9:       * 
    "00000010",  -- A:       * 
    "00000010",  -- B:       * 
    "11111100",  -- C: ******  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x3A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00011000",  -- 9:    **   
    "00011000",  -- A:    **   
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x3B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00011000",  -- 4:    **   
    "00011000",  -- 5:    **   
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00010000",  -- B:    *    
    "00100000",  -- C:   *     
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x3C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000010",  -- 4:       * 
    "00001100",  -- 5:     **  
    "00110000",  -- 6:   **    
    "11000000",  -- 7: **      
    "00110000",  -- 8:   **    
    "00001100",  -- 9:     **  
    "00000010",  -- A:       * 
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x3D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "11111110",  -- 4: ******* 
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "11111110",  -- A: ******* 
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x3E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "10000000",  -- 4: *       
    "01100000",  -- 5:  **     
    "00011000",  -- 6:    **   
    "00000110",  -- 7:      ** 
    "00011000",  -- 8:    **   
    "01100000",  -- 9:  **     
    "10000000",  -- A: *       
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x3F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111000",  -- 2:   ***   
    "01000100",  -- 3:  *   *  
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "00000010",  -- 6:       * 
    "00000100",  -- 7:      *  
    "00001000",  -- 8:     *   
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00000000",  -- B:         
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x40
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111000",  -- 2:   ***   
    "01000100",  -- 3:  *   *  
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10011110",  -- 6: *  **** 
    "10100010",  -- 7: * *   * 
    "10100010",  -- 8: * *   * 
    "10011110",  -- 9: *  **** 
    "10000000",  -- A: *       
    "01000010",  -- B:  *    * 
    "00111100",  -- C:   ****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x41
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00101000",  -- 3:   * *   
    "00101000",  -- 4:   * *   
    "00101000",  -- 5:   * *   
    "01000100",  -- 6:  *   *  
    "01111100",  -- 7:  *****  
    "01000100",  -- 8:  *   *  
    "01000100",  -- 9:  *   *  
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x42
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111100",  -- 2: ******  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000100",  -- 6: *    *  
    "11111000",  -- 7: *****   
    "10000100",  -- 8: *    *  
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "11111100",  -- C: ******  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x43
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "10000000",  -- 7: *       
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x44
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11110000",  -- 2: ****    
    "10001000",  -- 3: *   *   
    "10000100",  -- 4: *    *  
    "10000100",  -- 5: *    *  
    "10000010",  -- 6: *     * 
    "10000010",  -- 7: *     * 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000100",  -- A: *    *  
    "10000100",  -- B: *    *  
    "11111000",  -- C: *****   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x45
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111110",  -- 2: ******* 
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "11111100",  -- 7: ******  
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "11111110",  -- C: ******* 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x46
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111110",  -- 2: ******* 
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "11111100",  -- 7: ******  
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "10000000",  -- C: *       
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x47
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "10011110",  -- 7: *  **** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x48
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "01111100",  -- 7:  *****  
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x49
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111000",  -- 2:   ***   
    "00010000",  -- 3:    *    
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x4A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00011100",  -- 2:    ***  
    "00001000",  -- 3:     *   
    "00001000",  -- 4:     *   
    "00001000",  -- 5:     *   
    "00001000",  -- 6:     *   
    "00001000",  -- 7:     *   
    "00001000",  -- 8:     *   
    "00001000",  -- 9:     *   
    "10001000",  -- A: *   *   
    "10001000",  -- B: *   *   
    "01110000",  -- C:  ***    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x4B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "10000100",  -- 4: *    *  
    "10000100",  -- 5: *    *  
    "10001000",  -- 6: *   *   
    "11110000",  -- 7: ****    
    "10001000",  -- 8: *   *   
    "10000100",  -- 9: *    *  
    "10000100",  -- A: *    *  
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x4C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000000",  -- 2: *       
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "10000000",  -- 7: *       
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "11111110",  -- C: ******* 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x4D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "11000110",  -- 3: **   ** 
    "10101010",  -- 4: * * * * 
    "10101010",  -- 5: * * * * 
    "10101010",  -- 6: * * * * 
    "10010010",  -- 7: *  *  * 
    "10010010",  -- 8: *  *  * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x4E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "11000010",  -- 3: **    * 
    "10100010",  -- 4: * *   * 
    "10100010",  -- 5: * *   * 
    "10100010",  -- 6: * *   * 
    "10010010",  -- 7: *  *  * 
    "10001010",  -- 8: *   * * 
    "10001010",  -- 9: *   * * 
    "10001010",  -- A: *   * * 
    "10000110",  -- B: *    ** 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x4F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "10000010",  -- 7: *     * 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x50
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "11111100",  -- 7: ******  
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "10000000",  -- C: *       
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x51
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "10000010",  -- 7: *     * 
    "10000010",  -- 8: *     * 
    "10110010",  -- 9: * **  * 
    "10001010",  -- A: *   * * 
    "10000100",  -- B: *    *  
    "01111010",  -- C:  **** * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x52
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "11111100",  -- 7: ******  
    "10100000",  -- 8: * *     
    "10010000",  -- 9: *  *    
    "10001000",  -- A: *   *   
    "10000100",  -- B: *    *  
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x53
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "01111100",  -- 2:  *****  
    "10000010",  -- 3: *     * 
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000000",  -- 6: *       
    "01111100",  -- 7:  *****  
    "00000010",  -- 8:       * 
    "00000010",  -- 9:       * 
    "00000010",  -- A:       * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x54
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111110",  -- 2: ******* 
    "10010010",  -- 3: *  *  * 
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x55
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10000010",  -- 6: *     * 
    "10000010",  -- 7: *     * 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x56
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "01000100",  -- 5:  *   *  
    "01000100",  -- 6:  *   *  
    "01000100",  -- 7:  *   *  
    "00101000",  -- 8:   * *   
    "00101000",  -- 9:   * *   
    "00101000",  -- A:   * *   
    "00010000",  -- B:    *    
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x57
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "10000010",  -- 4: *     * 
    "10000010",  -- 5: *     * 
    "10010010",  -- 6: *  *  * 
    "10010010",  -- 7: *  *  * 
    "10101010",  -- 8: * * * * 
    "10101010",  -- 9: * * * * 
    "10101010",  -- A: * * * * 
    "11000110",  -- B: **   ** 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x58
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "01000100",  -- 4:  *   *  
    "01000100",  -- 5:  *   *  
    "00101000",  -- 6:   * *   
    "00111000",  -- 7:   ***   
    "00101000",  -- 8:   * *   
    "01000100",  -- 9:  *   *  
    "01000100",  -- A:  *   *  
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x59
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000010",  -- 2: *     * 
    "10000010",  -- 3: *     * 
    "01000100",  -- 4:  *   *  
    "01000100",  -- 5:  *   *  
    "00101000",  -- 6:   * *   
    "00101000",  -- 7:   * *   
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x5A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "11111110",  -- 2: ******* 
    "10000010",  -- 3: *     * 
    "00000100",  -- 4:      *  
    "00000100",  -- 5:      *  
    "00001000",  -- 6:     *   
    "00111000",  -- 7:   ***   
    "00100000",  -- 8:   *     
    "01000000",  -- 9:  *      
    "01000000",  -- A:  *      
    "10000010",  -- B: *     * 
    "11111110",  -- C: ******* 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x5B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111000",  -- 2:   ***   
    "00100000",  -- 3:   *     
    "00100000",  -- 4:   *     
    "00100000",  -- 5:   *     
    "00100000",  -- 6:   *     
    "00100000",  -- 7:   *     
    "00100000",  -- 8:   *     
    "00100000",  -- 9:   *     
    "00100000",  -- A:   *     
    "00100000",  -- B:   *     
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x5C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "10000000",  -- 4: *       
    "01000000",  -- 5:  *      
    "00100000",  -- 6:   *     
    "00010000",  -- 7:    *    
    "00001000",  -- 8:     *   
    "00000100",  -- 9:      *  
    "00000010",  -- A:       * 
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x5D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111000",  -- 2:   ***   
    "00001000",  -- 3:     *   
    "00001000",  -- 4:     *   
    "00001000",  -- 5:     *   
    "00001000",  -- 6:     *   
    "00001000",  -- 7:     *   
    "00001000",  -- 8:     *   
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00001000",  -- B:     *   
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x5E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00010000",  -- 3:    *    
    "00101000",  -- 4:   * *   
    "01000100",  -- 5:  *   *  
    "10000010",  -- 6: *     * 
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x5F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "11111110",  -- C: ******* 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x60
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00100000",  -- 2:   *     
    "00100000",  -- 3:   *     
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00001000",  -- 6:     *   
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x61
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00111010",  -- 6:   *** * 
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "11000110",  -- B: **   ** 
    "00111010",  -- C:   *** * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x62
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000000",  -- 2: *       
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10111000",  -- 6: * ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "11000110",  -- B: **   ** 
    "10111000",  -- C: * ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x63
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00111100",  -- 6:   ****  
    "11000010",  -- 7: **    * 
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "11000010",  -- B: **    * 
    "00111100",  -- C:   ****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x64
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000010",  -- 2:       * 
    "00000010",  -- 3:       * 
    "00000010",  -- 4:       * 
    "00000010",  -- 5:       * 
    "00111010",  -- 6:   *** * 
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "11000110",  -- B: **   ** 
    "00111010",  -- C:   *** * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x65
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00111000",  -- 6:   ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "11111100",  -- 9: ******  
    "10000000",  -- A: *       
    "11000110",  -- B: **   ** 
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x66
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00111100",  -- 2:   ****  
    "01000010",  -- 3:  *    * 
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "11111000",  -- 6: *****   
    "10000000",  -- 7: *       
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "10000000",  -- C: *       
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x67
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00111000",  -- 6:   ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "01111110",  -- 9:  ****** 
    "00000010",  -- A:       * 
    "11000110",  -- B: **   ** 
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x68
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000000",  -- 2: *       
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10111000",  -- 6: * ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x69
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00010000",  -- 3:    *    
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00010000",  -- 6:    *    
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010010",  -- B:    *  * 
    "00001100",  -- C:     **  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x6A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000100",  -- 3:      *  
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000100",  -- 6:      *  
    "00000100",  -- 7:      *  
    "00000100",  -- 8:      *  
    "00000100",  -- 9:      *  
    "00000100",  -- A:      *  
    "10001000",  -- B: *   *   
    "01110000",  -- C:  ***    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x6B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "10000110",  -- 6: *    ** 
    "10111000",  -- 7: * ***   
    "11000000",  -- 8: **      
    "10110000",  -- 9: * **    
    "10001000",  -- A: *   *   
    "10000100",  -- B: *    *  
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x6C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00100000",  -- 2:   *     
    "00100000",  -- 3:   *     
    "00100000",  -- 4:   *     
    "00100000",  -- 5:   *     
    "00100000",  -- 6:   *     
    "00100000",  -- 7:   *     
    "00100000",  -- 8:   *     
    "00100000",  -- 9:   *     
    "00100000",  -- A:   *     
    "00010000",  -- B:    *    
    "00001110",  -- C:     *** 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x6D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10101100",  -- 6: * * **  
    "11010010",  -- 7: ** *  * 
    "10010010",  -- 8: *  *  * 
    "10010010",  -- 9: *  *  * 
    "10010010",  -- A: *  *  * 
    "10010010",  -- B: *  *  * 
    "10010010",  -- C: *  *  * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x6E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10111000",  -- 6: * ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "10000010",  -- B: *     * 
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x6F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00111000",  -- 6:   ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "11000110",  -- B: **   ** 
    "00111000",  -- C:   ***   
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x70
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10111000",  -- 6: * ***   
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "11111100",  -- 9: ******  
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "10000000",  -- C: *       
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x71
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00111010",  -- 6:   *** * 
    "11000110",  -- 7: **   ** 
    "10000010",  -- 8: *     * 
    "01111110",  -- 9:  ****** 
    "00000010",  -- A:       * 
    "00000010",  -- B:       * 
    "00000010",  -- C:       * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x72
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10111000",  -- 6: * ***   
    "11000110",  -- 7: **   ** 
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "10000000",  -- B: *       
    "10000000",  -- C: *       
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x73
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "01111100",  -- 6:  *****  
    "10000010",  -- 7: *     * 
    "10000000",  -- 8: *       
    "01111110",  -- 9:  ****** 
    "00000010",  -- A:       * 
    "10000010",  -- B: *     * 
    "01111100",  -- C:  *****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x74
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "10000000",  -- 2: *       
    "10000000",  -- 3: *       
    "10000000",  -- 4: *       
    "10000000",  -- 5: *       
    "11111000",  -- 6: *****   
    "10000000",  -- 7: *       
    "10000000",  -- 8: *       
    "10000000",  -- 9: *       
    "10000000",  -- A: *       
    "01000010",  -- B:  *    * 
    "00111100",  -- C:   ****  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x75
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10000010",  -- 6: *     * 
    "10000010",  -- 7: *     * 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "10000010",  -- A: *     * 
    "11000110",  -- B: **   ** 
    "00111010",  -- C:   *** * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x76
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10000010",  -- 6: *     * 
    "10000010",  -- 7: *     * 
    "10000010",  -- 8: *     * 
    "10000010",  -- 9: *     * 
    "01000100",  -- A:  *   *  
    "00101000",  -- B:   * *   
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x77
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "10000010",  -- 6: *     * 
    "10010010",  -- 7: *  *  * 
    "10010010",  -- 8: *  *  * 
    "10010010",  -- 9: *  *  * 
    "10010010",  -- A: *  *  * 
    "10010010",  -- B: *  *  * 
    "01101100",  -- C:  ** **  
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x78
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "10000010",  -- 7: *     * 
    "01000100",  -- 8:  *   *  
    "00101000",  -- 9:   * *   
    "00111000",  -- A:   ***   
    "01000100",  -- B:  *   *  
    "10000010",  -- C: *     * 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x79
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "10000010",  -- 7: *     * 
    "01000010",  -- 8:  *    * 
    "00111100",  -- 9:   ****  
    "00001000",  -- A:     *   
    "00001000",  -- B:     *   
    "00110000",  -- C:   **    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x7A
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "11111110",  -- 7: ******* 
    "00000100",  -- 8:      *  
    "00001000",  -- 9:     *   
    "00110000",  -- A:   **    
    "01000000",  -- B:  *      
    "11111110",  -- C: ******* 
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x7B
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00100000",  -- 3:   *     
    "00100000",  -- 4:   *     
    "00100000",  -- 5:   *     
    "01000000",  -- 6:  *      
    "10000000",  -- 7: *       
    "01000000",  -- 8:  *      
    "00100000",  -- 9:   *     
    "00100000",  -- A:   *     
    "00100000",  -- B:   *     
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x7C
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00010000",  -- 3:    *    
    "00010000",  -- 4:    *    
    "00010000",  -- 5:    *    
    "00010000",  -- 6:    *    
    "00010000",  -- 7:    *    
    "00010000",  -- 8:    *    
    "00010000",  -- 9:    *    
    "00010000",  -- A:    *    
    "00010000",  -- B:    *    
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x7D
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00010000",  -- 2:    *    
    "00001000",  -- 3:     *   
    "00001000",  -- 4:     *   
    "00001000",  -- 5:     *   
    "00000100",  -- 6:      *  
    "00000010",  -- 7:       * 
    "00000100",  -- 8:      *  
    "00001000",  -- 9:     *   
    "00001000",  -- A:     *   
    "00001000",  -- B:     *   
    "00010000",  -- C:    *    
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x7E
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "01100000",  -- 6:  **     
    "10010010",  -- 7: *  *  * 
    "00001100",  -- 8:     **  
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
      -- Char Code: 0x7F
    "00000000",  -- 0:         
    "00000000",  -- 1:         
    "00000000",  -- 2:         
    "00000000",  -- 3:         
    "00000000",  -- 4:         
    "00000000",  -- 5:         
    "00000000",  -- 6:         
    "00000000",  -- 7:         
    "00000000",  -- 8:         
    "00000000",  -- 9:         
    "00000000",  -- A:         
    "00000000",  -- B:         
    "00000000",  -- C:         
    "00000000",  -- D:         
    "00000000",  -- E:         
    "00000000",  -- F:         
    others => "00000000"
  );

  constant FONT_8X16X128_2 : Font_type := (
    ID       => 3,
    Width    => 8,
    Height   => 16,
    NumChars => 128,
    Data     => FONT_ROM_8X16X128_2
  );
  
-- More font tables to be added later?
  
end font_pack;


package body font_pack is

end font_pack;
